

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n449) );
  XNOR2_X1 U324 ( .A(n450), .B(n449), .ZN(n457) );
  NOR2_X1 U325 ( .A1(n451), .A2(n403), .ZN(n404) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n520) );
  XOR2_X1 U327 ( .A(G211GAT), .B(KEYINPUT21), .Z(n291) );
  XOR2_X1 U328 ( .A(n363), .B(n362), .Z(n292) );
  XNOR2_X1 U329 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U330 ( .A(n430), .B(n429), .ZN(n434) );
  NOR2_X1 U331 ( .A1(n535), .A2(n492), .ZN(n521) );
  XNOR2_X1 U332 ( .A(n373), .B(n372), .ZN(n374) );
  NOR2_X1 U333 ( .A1(n461), .A2(n460), .ZN(n566) );
  XOR2_X1 U334 ( .A(n458), .B(KEYINPUT48), .Z(n536) );
  XNOR2_X1 U335 ( .A(n375), .B(n374), .ZN(n391) );
  XOR2_X1 U336 ( .A(KEYINPUT38), .B(n439), .Z(n493) );
  XNOR2_X1 U337 ( .A(n465), .B(G183GAT), .ZN(n466) );
  XNOR2_X1 U338 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U339 ( .A(n467), .B(n466), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n443), .B(n442), .ZN(G1328GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT5), .B(G57GAT), .Z(n294) );
  XNOR2_X1 U342 ( .A(KEYINPUT88), .B(KEYINPUT6), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n300) );
  XOR2_X1 U344 ( .A(G155GAT), .B(KEYINPUT2), .Z(n296) );
  XNOR2_X1 U345 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n365) );
  XOR2_X1 U347 ( .A(G85GAT), .B(n365), .Z(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT0), .B(G127GAT), .Z(n379) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(n379), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n313) );
  XOR2_X1 U352 ( .A(G162GAT), .B(G120GAT), .Z(n302) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G113GAT), .ZN(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U355 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n304) );
  XNOR2_X1 U356 ( .A(G1GAT), .B(G148GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U359 ( .A(KEYINPUT85), .B(KEYINPUT4), .Z(n308) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U362 ( .A(KEYINPUT1), .B(n309), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n461) );
  XOR2_X1 U365 ( .A(G50GAT), .B(G162GAT), .Z(n363) );
  XNOR2_X1 U366 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n314), .B(KEYINPUT7), .ZN(n410) );
  XOR2_X1 U368 ( .A(n363), .B(n410), .Z(n316) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n317), .B(KEYINPUT9), .ZN(n319) );
  XOR2_X1 U372 ( .A(G36GAT), .B(G218GAT), .Z(n358) );
  XOR2_X1 U373 ( .A(n358), .B(KEYINPUT11), .Z(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n321) );
  XNOR2_X1 U376 ( .A(KEYINPUT10), .B(KEYINPUT72), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n328) );
  XNOR2_X1 U379 ( .A(G43GAT), .B(G190GAT), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n324), .B(G134GAT), .ZN(n380) );
  XOR2_X1 U381 ( .A(G92GAT), .B(G85GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n424) );
  XNOR2_X1 U384 ( .A(n380), .B(n424), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n548) );
  XNOR2_X1 U386 ( .A(n548), .B(KEYINPUT73), .ZN(n559) );
  XNOR2_X1 U387 ( .A(KEYINPUT36), .B(n559), .ZN(n451) );
  XOR2_X1 U388 ( .A(G57GAT), .B(KEYINPUT13), .Z(n428) );
  XOR2_X1 U389 ( .A(G71GAT), .B(G127GAT), .Z(n330) );
  XNOR2_X1 U390 ( .A(G15GAT), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U392 ( .A(n428), .B(n331), .Z(n333) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n334), .B(KEYINPUT75), .Z(n337) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G1GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n335), .B(G8GAT), .ZN(n407) );
  XNOR2_X1 U398 ( .A(n407), .B(KEYINPUT74), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n345) );
  XOR2_X1 U400 ( .A(G64GAT), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U401 ( .A(G78GAT), .B(G155GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n341) );
  XNOR2_X1 U404 ( .A(KEYINPUT12), .B(KEYINPUT76), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U406 ( .A(n343), .B(n342), .Z(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n577) );
  XOR2_X1 U408 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n347) );
  XNOR2_X1 U409 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U411 ( .A(n348), .B(G183GAT), .Z(n350) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G176GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n388) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(KEYINPUT84), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n291), .B(n351), .ZN(n362) );
  XOR2_X1 U416 ( .A(n362), .B(G8GAT), .Z(n353) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U419 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n355) );
  XNOR2_X1 U420 ( .A(G190GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U422 ( .A(n357), .B(n356), .Z(n360) );
  XOR2_X1 U423 ( .A(G204GAT), .B(G64GAT), .Z(n435) );
  XNOR2_X1 U424 ( .A(n358), .B(n435), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n388), .B(n361), .ZN(n512) );
  XOR2_X1 U427 ( .A(KEYINPUT27), .B(n512), .Z(n397) );
  NAND2_X1 U428 ( .A1(n461), .A2(n397), .ZN(n535) );
  NAND2_X1 U429 ( .A1(G228GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n292), .B(n364), .ZN(n366) );
  XOR2_X1 U431 ( .A(n366), .B(n365), .Z(n368) );
  XNOR2_X1 U432 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U434 ( .A(G148GAT), .B(G78GAT), .Z(n436) );
  XOR2_X1 U435 ( .A(n369), .B(n436), .Z(n375) );
  XOR2_X1 U436 ( .A(KEYINPUT24), .B(G204GAT), .Z(n371) );
  XNOR2_X1 U437 ( .A(KEYINPUT23), .B(KEYINPUT83), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n373) );
  XNOR2_X1 U439 ( .A(G218GAT), .B(G106GAT), .ZN(n372) );
  XOR2_X1 U440 ( .A(KEYINPUT28), .B(n391), .Z(n492) );
  XOR2_X1 U441 ( .A(n521), .B(KEYINPUT91), .Z(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT79), .B(KEYINPUT20), .Z(n377) );
  NAND2_X1 U443 ( .A1(G227GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U445 ( .A(KEYINPUT81), .B(n378), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U447 ( .A(G120GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U448 ( .A(n381), .B(n423), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U450 ( .A(n384), .B(KEYINPUT78), .Z(n386) );
  XOR2_X1 U451 ( .A(G113GAT), .B(G15GAT), .Z(n406) );
  XNOR2_X1 U452 ( .A(n406), .B(G99GAT), .ZN(n385) );
  XNOR2_X1 U453 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U454 ( .A(KEYINPUT82), .B(n520), .Z(n389) );
  NAND2_X1 U455 ( .A1(n390), .A2(n389), .ZN(n402) );
  INV_X1 U456 ( .A(n512), .ZN(n485) );
  NAND2_X1 U457 ( .A1(n520), .A2(n485), .ZN(n392) );
  NAND2_X1 U458 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n393), .B(KEYINPUT93), .ZN(n394) );
  XNOR2_X1 U460 ( .A(KEYINPUT25), .B(n394), .ZN(n399) );
  NOR2_X1 U461 ( .A1(n520), .A2(n391), .ZN(n396) );
  XNOR2_X1 U462 ( .A(KEYINPUT92), .B(KEYINPUT26), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n565) );
  NAND2_X1 U464 ( .A1(n397), .A2(n565), .ZN(n398) );
  NAND2_X1 U465 ( .A1(n399), .A2(n398), .ZN(n400) );
  INV_X1 U466 ( .A(n461), .ZN(n509) );
  NAND2_X1 U467 ( .A1(n400), .A2(n509), .ZN(n401) );
  NAND2_X1 U468 ( .A1(n402), .A2(n401), .ZN(n471) );
  NAND2_X1 U469 ( .A1(n577), .A2(n471), .ZN(n403) );
  XOR2_X1 U470 ( .A(KEYINPUT100), .B(n404), .Z(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT37), .B(n405), .ZN(n507) );
  XOR2_X1 U472 ( .A(n407), .B(n406), .Z(n409) );
  XNOR2_X1 U473 ( .A(G43GAT), .B(G50GAT), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U475 ( .A(n410), .B(KEYINPUT66), .Z(n412) );
  NAND2_X1 U476 ( .A1(G229GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U478 ( .A(n414), .B(n413), .Z(n422) );
  XOR2_X1 U479 ( .A(G197GAT), .B(G141GAT), .Z(n416) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G36GAT), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n418) );
  XNOR2_X1 U483 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n567) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n426) );
  NAND2_X1 U488 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U490 ( .A(G176GAT), .B(KEYINPUT31), .ZN(n427) );
  XOR2_X1 U491 ( .A(KEYINPUT32), .B(KEYINPUT68), .Z(n432) );
  XNOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n431) );
  XOR2_X1 U493 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n444) );
  INV_X1 U497 ( .A(n444), .ZN(n572) );
  NOR2_X1 U498 ( .A1(n567), .A2(n444), .ZN(n472) );
  NAND2_X1 U499 ( .A1(n507), .A2(n472), .ZN(n439) );
  NAND2_X1 U500 ( .A1(n461), .A2(n493), .ZN(n443) );
  XOR2_X1 U501 ( .A(G29GAT), .B(KEYINPUT99), .Z(n441) );
  XNOR2_X1 U502 ( .A(KEYINPUT101), .B(KEYINPUT39), .ZN(n440) );
  INV_X1 U503 ( .A(n567), .ZN(n523) );
  XOR2_X1 U504 ( .A(KEYINPUT41), .B(n444), .Z(n525) );
  AND2_X1 U505 ( .A1(n523), .A2(n525), .ZN(n446) );
  XNOR2_X1 U506 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U508 ( .A(n577), .ZN(n528) );
  OR2_X1 U509 ( .A1(n548), .A2(n528), .ZN(n447) );
  OR2_X1 U510 ( .A1(n448), .A2(n447), .ZN(n450) );
  XOR2_X1 U511 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n453) );
  NOR2_X1 U512 ( .A1(n577), .A2(n451), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U514 ( .A1(n454), .A2(n444), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n455), .A2(n567), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n457), .A2(n456), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n512), .A2(n536), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT54), .B(n459), .Z(n460) );
  NAND2_X1 U519 ( .A1(n566), .A2(n391), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n462) );
  XNOR2_X1 U521 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n464), .A2(n520), .ZN(n558) );
  NOR2_X1 U523 ( .A1(n577), .A2(n558), .ZN(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n465) );
  INV_X1 U525 ( .A(n559), .ZN(n531) );
  NOR2_X1 U526 ( .A1(n577), .A2(n531), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT77), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n469), .Z(n470) );
  AND2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n496) );
  NAND2_X1 U530 ( .A1(n472), .A2(n496), .ZN(n481) );
  NOR2_X1 U531 ( .A1(n509), .A2(n481), .ZN(n474) );
  XNOR2_X1 U532 ( .A(KEYINPUT34), .B(KEYINPUT94), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U535 ( .A1(n512), .A2(n481), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n476) );
  XNOR2_X1 U537 ( .A(n477), .B(n476), .ZN(G1325GAT) );
  INV_X1 U538 ( .A(n520), .ZN(n514) );
  NOR2_X1 U539 ( .A1(n514), .A2(n481), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT96), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  INV_X1 U543 ( .A(n492), .ZN(n517) );
  NOR2_X1 U544 ( .A1(n517), .A2(n481), .ZN(n483) );
  XNOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NAND2_X1 U548 ( .A1(n493), .A2(n485), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n486), .B(KEYINPUT102), .ZN(n487) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n487), .ZN(G1329GAT) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(KEYINPUT103), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n489) );
  NAND2_X1 U553 ( .A1(n493), .A2(n520), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n525), .ZN(n555) );
  NOR2_X1 U560 ( .A1(n523), .A2(n555), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n508), .A2(n496), .ZN(n503) );
  NOR2_X1 U562 ( .A1(n509), .A2(n503), .ZN(n498) );
  XNOR2_X1 U563 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U564 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n499), .Z(G1332GAT) );
  NOR2_X1 U566 ( .A1(n512), .A2(n503), .ZN(n500) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n500), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n514), .A2(n503), .ZN(n502) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(KEYINPUT107), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n517), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(KEYINPUT43), .B(KEYINPUT108), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n506), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n516) );
  NOR2_X1 U576 ( .A1(n509), .A2(n516), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n512), .A2(n516), .ZN(n513) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n513), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U587 ( .A1(n536), .A2(n522), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n523), .A2(n532), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U591 ( .A1(n532), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  NAND2_X1 U593 ( .A1(n532), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n565), .A2(n537), .ZN(n547) );
  NOR2_X1 U601 ( .A1(n567), .A2(n547), .ZN(n538) );
  XOR2_X1 U602 ( .A(G141GAT), .B(n538), .Z(G1344GAT) );
  NOR2_X1 U603 ( .A1(n555), .A2(n547), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT113), .Z(n540) );
  XNOR2_X1 U605 ( .A(G148GAT), .B(KEYINPUT112), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT52), .B(n541), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n577), .A2(n547), .ZN(n545) );
  XNOR2_X1 U610 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n546), .ZN(G1346GAT) );
  INV_X1 U613 ( .A(n547), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(KEYINPUT116), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n551), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n567), .A2(n558), .ZN(n552) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n554) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n555), .A2(n558), .ZN(n556) );
  XOR2_X1 U623 ( .A(n557), .B(n556), .Z(G1349GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n564) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n561) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT121), .B(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1351GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT124), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n580) );
  NOR2_X1 U632 ( .A1(n567), .A2(n580), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n580), .A2(n572), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n574) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n580), .ZN(n579) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n451), .A2(n580), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

