//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G57gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT97), .ZN(new_n204));
  INV_X1    g003(.A(G57gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G64gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT98), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(KEYINPUT97), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(KEYINPUT98), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n204), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G71gat), .B(G78gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT99), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n203), .B2(new_n206), .ZN(new_n217));
  NOR2_X1   g016(.A1(G71gat), .A2(G78gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT96), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(new_n213), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n220), .C1(new_n219), .C2(new_n213), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G231gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(G127gat), .B(G155gat), .Z(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT100), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n226), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G1gat), .B2(new_n230), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n222), .B2(new_n223), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT101), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n229), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n239));
  XNOR2_X1  g038(.A(G183gat), .B(G211gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n238), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G43gat), .B(G50gat), .Z(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT92), .Z(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT90), .B(KEYINPUT14), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  INV_X1    g048(.A(G36gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n252));
  AOI211_X1 g051(.A(G29gat), .B(G36gat), .C1(new_n252), .C2(KEYINPUT14), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n244), .A2(new_n245), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(G29gat), .B2(G36gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n247), .A2(KEYINPUT93), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT93), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n256), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n246), .B(KEYINPUT92), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT91), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n254), .A2(new_n263), .B1(G29gat), .B2(G36gat), .ZN(new_n264));
  OR3_X1    g063(.A1(new_n251), .A2(new_n263), .A3(new_n253), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n261), .A2(new_n257), .B1(new_n266), .B2(new_n255), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT17), .ZN(new_n272));
  NAND2_X1  g071(.A1(G85gat), .A2(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT7), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  INV_X1    g074(.A(G85gat), .ZN(new_n276));
  INV_X1    g075(.A(G92gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(KEYINPUT8), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G99gat), .B(G106gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND3_X1  g080(.A1(new_n270), .A2(new_n272), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  AND2_X1   g082(.A1(G232gat), .A2(G233gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n268), .A2(new_n283), .B1(KEYINPUT41), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT103), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n286), .B(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n284), .A2(KEYINPUT41), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT102), .ZN(new_n292));
  XNOR2_X1  g091(.A(G134gat), .B(G162gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n290), .B(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n281), .B(new_n222), .Z(new_n296));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n216), .A4(new_n221), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n296), .A2(new_n301), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT104), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n302), .A2(KEYINPUT104), .A3(new_n304), .A4(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n307), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n298), .A2(new_n299), .B1(G230gat), .B2(G233gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n303), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n243), .A2(new_n295), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G229gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n235), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n268), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n235), .B1(new_n271), .B2(KEYINPUT17), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n268), .A2(new_n269), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n319), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT18), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT94), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n320), .B1(new_n268), .B2(new_n269), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n327), .A2(new_n272), .B1(new_n268), .B2(new_n320), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT94), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT18), .A4(new_n319), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n271), .A2(new_n235), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n321), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n319), .B(KEYINPUT13), .Z(new_n334));
  AOI22_X1  g133(.A1(new_n324), .A2(new_n325), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G113gat), .B(G141gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n337), .B(G197gat), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT11), .B(G169gat), .Z(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n340), .B(KEYINPUT12), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n331), .A2(new_n335), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT72), .ZN(new_n347));
  INV_X1    g146(.A(G211gat), .ZN(new_n348));
  INV_X1    g147(.A(G218gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT71), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT71), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G218gat), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n348), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n347), .B1(new_n353), .B2(KEYINPUT22), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT22), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT71), .B(G218gat), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT72), .B(new_n355), .C1(new_n356), .C2(new_n348), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(G197gat), .B(G204gat), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n346), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n346), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n359), .B(new_n362), .C1(new_n354), .C2(new_n357), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(G183gat), .A3(G190gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G183gat), .B(G190gat), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT64), .B(new_n368), .C1(new_n369), .C2(new_n367), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n368), .B1(new_n369), .B2(new_n367), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT23), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT24), .ZN(new_n381));
  INV_X1    g180(.A(G183gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n381), .B1(new_n386), .B2(KEYINPUT24), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n387), .B(new_n388), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(KEYINPUT27), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G183gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n393), .A3(new_n384), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT28), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT28), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n396), .A4(new_n384), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n395), .A2(new_n380), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n399));
  OR3_X1    g198(.A1(new_n399), .A2(new_n373), .A3(KEYINPUT65), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT65), .B1(new_n399), .B2(new_n373), .ZN(new_n401));
  INV_X1    g200(.A(new_n373), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n401), .C1(KEYINPUT26), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n390), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n406));
  AOI21_X1  g205(.A(new_n366), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n389), .A2(new_n379), .B1(new_n398), .B2(new_n403), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(new_n365), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n364), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n365), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n361), .A2(new_n363), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n405), .A2(new_n366), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n410), .A2(KEYINPUT75), .A3(new_n414), .A4(new_n417), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT76), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n420), .A2(KEYINPUT76), .A3(new_n421), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429));
  INV_X1    g228(.A(G141gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(G148gat), .ZN(new_n431));
  INV_X1    g230(.A(G148gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(G141gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G155gat), .B(G162gat), .Z(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G155gat), .ZN(new_n437));
  INV_X1    g236(.A(G162gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G141gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n443), .A3(G148gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n431), .ZN(new_n445));
  AOI221_X4 g244(.A(KEYINPUT78), .B1(new_n439), .B2(new_n440), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n445), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n440), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n436), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G113gat), .ZN(new_n452));
  INV_X1    g251(.A(G120gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n455));
  NAND2_X1  g254(.A1(G113gat), .A2(G120gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(G127gat), .A2(G134gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(G127gat), .A2(G134gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(G113gat), .A2(G120gat), .ZN(new_n462));
  NOR2_X1   g261(.A1(G113gat), .A2(G120gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT67), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n465), .A3(new_n456), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n466), .A3(new_n455), .ZN(new_n467));
  INV_X1    g266(.A(G127gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G127gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n459), .B1(new_n472), .B2(G134gat), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n461), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n474), .B(new_n436), .C1(new_n450), .C2(new_n446), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n428), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT77), .B(G141gat), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n431), .B1(new_n483), .B2(G148gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n449), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT78), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n448), .A2(new_n447), .A3(new_n449), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n486), .A2(new_n487), .B1(new_n434), .B2(new_n435), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n475), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n451), .A2(KEYINPUT3), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n482), .B(new_n479), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT79), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n487), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n436), .A4(new_n474), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n481), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n488), .A2(new_n489), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n451), .A2(KEYINPUT3), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n475), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n497), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n428), .A4(new_n479), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G1gat), .B(G29gat), .Z(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G57gat), .B(G85gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g311(.A(new_n510), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n499), .A2(new_n513), .A3(new_n504), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n510), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n410), .A2(new_n414), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(KEYINPUT74), .A3(KEYINPUT30), .A4(new_n417), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n418), .B2(new_n421), .ZN(new_n521));
  INV_X1    g320(.A(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(new_n417), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n519), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n427), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT35), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n408), .B(new_n474), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(G227gat), .B2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT34), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(G227gat), .A3(G233gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n534));
  XOR2_X1   g333(.A(G71gat), .B(G99gat), .Z(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G43gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n533), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT68), .B(KEYINPUT33), .Z(new_n539));
  OAI211_X1 g338(.A(new_n534), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(new_n541), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n545), .A3(new_n540), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT83), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n412), .B1(new_n500), .B2(new_n406), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n406), .B1(new_n361), .B2(new_n363), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT82), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(new_n406), .C1(new_n361), .C2(new_n363), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n489), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n556), .B2(new_n451), .ZN(new_n557));
  INV_X1    g356(.A(G228gat), .ZN(new_n558));
  INV_X1    g357(.A(G233gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n550), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT3), .B1(new_n552), .B2(KEYINPUT82), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n488), .B1(new_n563), .B2(new_n555), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT83), .B(new_n562), .C1(new_n564), .C2(new_n551), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n500), .A2(new_n406), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n560), .B1(new_n567), .B2(new_n412), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n364), .A2(new_n569), .A3(KEYINPUT29), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n489), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(new_n572), .B2(new_n451), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n566), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G22gat), .ZN(new_n576));
  INV_X1    g375(.A(G22gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n566), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G78gat), .B(G106gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G50gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n576), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n582), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n577), .B1(new_n566), .B2(new_n574), .ZN(new_n585));
  AOI211_X1 g384(.A(G22gat), .B(new_n573), .C1(new_n561), .C2(new_n565), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n549), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n528), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n591));
  AOI211_X1 g390(.A(new_n549), .B(new_n525), .C1(new_n583), .C2(new_n587), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n549), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n582), .B1(new_n576), .B2(new_n578), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n585), .A2(new_n586), .A3(new_n584), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n526), .B(new_n595), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT89), .A3(KEYINPUT35), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n590), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n502), .A2(new_n503), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n480), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT39), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n602), .B(KEYINPUT39), .C1(new_n480), .C2(new_n478), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT85), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT40), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n603), .A2(new_n604), .A3(new_n513), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n511), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n604), .A3(new_n513), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n427), .A2(new_n524), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n523), .A2(KEYINPUT37), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n518), .B2(new_n417), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618));
  INV_X1    g417(.A(new_n407), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n364), .B1(new_n619), .B2(new_n413), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n411), .A2(new_n364), .A3(new_n413), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT37), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n618), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n420), .B(new_n422), .C1(new_n617), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n522), .A2(KEYINPUT37), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n618), .B1(new_n625), .B2(new_n616), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT87), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n517), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n583), .A2(new_n587), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT86), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n612), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n614), .A2(new_n631), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT70), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n549), .A2(new_n637), .A3(KEYINPUT36), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT36), .B1(new_n549), .B2(new_n637), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n583), .A2(new_n587), .A3(new_n525), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n345), .B1(new_n600), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT95), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n528), .A2(new_n588), .A3(new_n589), .ZN(new_n646));
  AOI211_X1 g445(.A(new_n591), .B(new_n593), .C1(new_n588), .C2(new_n526), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT89), .B1(new_n598), .B2(KEYINPUT35), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n635), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n345), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n318), .B1(new_n645), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n629), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n645), .A2(new_n654), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  AND4_X1   g459(.A1(new_n612), .A2(new_n659), .A3(new_n317), .A4(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n234), .B1(new_n655), .B2(new_n612), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT42), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n659), .A2(new_n612), .A3(new_n317), .A4(new_n660), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n658), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n653), .B1(new_n652), .B2(new_n345), .ZN(new_n668));
  INV_X1    g467(.A(new_n345), .ZN(new_n669));
  AOI211_X1 g468(.A(KEYINPUT95), .B(new_n669), .C1(new_n649), .C2(new_n651), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n612), .B(new_n317), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(G8gat), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n665), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  INV_X1    g472(.A(new_n612), .ZN(new_n674));
  AOI211_X1 g473(.A(new_n674), .B(new_n318), .C1(new_n645), .C2(new_n654), .ZN(new_n675));
  AOI21_X1  g474(.A(KEYINPUT42), .B1(new_n675), .B2(new_n660), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n673), .A2(new_n676), .A3(KEYINPUT105), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n667), .A2(new_n677), .ZN(G1325gat));
  AOI21_X1  g477(.A(G15gat), .B1(new_n655), .B2(new_n595), .ZN(new_n679));
  INV_X1    g478(.A(new_n640), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT106), .Z(new_n682));
  AOI21_X1  g481(.A(new_n679), .B1(new_n655), .B2(new_n682), .ZN(G1326gat));
  INV_X1    g482(.A(new_n632), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n655), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  INV_X1    g486(.A(new_n295), .ZN(new_n688));
  INV_X1    g487(.A(new_n316), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n243), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n688), .B(new_n690), .C1(new_n645), .C2(new_n654), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n249), .A3(new_n629), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT107), .B1(new_n636), .B2(new_n642), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n650), .A2(new_n697), .A3(new_n635), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n649), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n699), .B2(new_n688), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n295), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n690), .A2(new_n669), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n517), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n692), .A2(new_n693), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n694), .A2(new_n704), .A3(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n250), .A3(new_n612), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n703), .B2(new_n674), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(KEYINPUT46), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n712), .A3(new_n595), .ZN(new_n713));
  OAI21_X1  g512(.A(G43gat), .B1(new_n703), .B2(new_n640), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1330gat));
  NOR2_X1   g516(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n632), .A2(G50gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n691), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G50gat), .B1(new_n703), .B2(new_n632), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1331gat));
  NAND4_X1  g523(.A1(new_n669), .A2(new_n688), .A3(new_n242), .A4(new_n316), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n699), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n629), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g527(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT49), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(new_n202), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n726), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n202), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1333gat));
  NAND2_X1  g537(.A1(new_n726), .A2(new_n595), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  AOI21_X1  g539(.A(G71gat), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n726), .A2(G71gat), .A3(new_n680), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT50), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1334gat));
  NAND2_X1  g547(.A1(new_n726), .A2(new_n684), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g549(.A1(new_n345), .A2(new_n242), .A3(new_n689), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n700), .A2(new_n701), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n517), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n649), .A2(new_n696), .A3(new_n698), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n345), .A2(new_n242), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n295), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n295), .A4(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n316), .A2(new_n276), .A3(new_n629), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n753), .B1(new_n761), .B2(new_n762), .ZN(G1336gat));
  NAND4_X1  g562(.A1(new_n700), .A2(new_n612), .A3(new_n701), .A4(new_n751), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n765), .A3(G92gat), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n764), .B2(G92gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n756), .A2(new_n768), .A3(KEYINPUT51), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT51), .B1(new_n756), .B2(new_n768), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n731), .A2(G92gat), .A3(new_n689), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n766), .A2(new_n767), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(G92gat), .B1(new_n752), .B2(new_n731), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(new_n760), .B2(new_n771), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(KEYINPUT114), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n776), .B2(new_n777), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n774), .A2(new_n775), .B1(new_n778), .B2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n752), .B2(new_n640), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n689), .A2(G99gat), .A3(new_n549), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n761), .B2(new_n782), .ZN(G1338gat));
  OAI21_X1  g582(.A(G106gat), .B1(new_n752), .B2(new_n632), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n632), .A2(new_n689), .A3(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n760), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n769), .A2(new_n770), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n785), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(new_n784), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n307), .B1(new_n314), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n302), .A2(KEYINPUT54), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n300), .A2(new_n301), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n794), .B(KEYINPUT55), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(new_n312), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n345), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n328), .A2(new_n319), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n333), .A2(new_n334), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n340), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n316), .A2(new_n344), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n295), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n344), .A2(new_n295), .A3(new_n801), .A4(new_n805), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n243), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n317), .A2(new_n669), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n811), .A2(new_n517), .A3(new_n684), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n732), .A2(new_n549), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n669), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(new_n452), .ZN(G1340gat));
  NOR2_X1   g615(.A1(new_n814), .A2(new_n689), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(new_n453), .ZN(G1341gat));
  NOR2_X1   g617(.A1(new_n814), .A2(new_n243), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n472), .A2(KEYINPUT115), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(G1342gat));
  NOR2_X1   g620(.A1(new_n688), .A2(new_n612), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  AOI211_X1 g622(.A(G134gat), .B(new_n549), .C1(new_n823), .C2(KEYINPUT56), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n812), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n825), .A2(new_n823), .A3(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n823), .B2(KEYINPUT56), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n295), .A3(new_n813), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n829), .B2(G134gat), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n829), .A2(new_n828), .A3(G134gat), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n826), .B(new_n827), .C1(new_n830), .C2(new_n831), .ZN(G1343gat));
  AOI21_X1  g631(.A(new_n632), .B1(new_n809), .B2(new_n810), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n680), .A2(new_n517), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n669), .A2(G141gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n833), .A2(new_n731), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT119), .Z(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n731), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n811), .B2(new_n632), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n316), .A2(new_n842), .A3(new_n344), .A4(new_n805), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n802), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n808), .B1(new_n844), .B2(new_n688), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n810), .B1(new_n845), .B2(new_n242), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n632), .A2(new_n839), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n838), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n483), .B1(new_n849), .B2(new_n345), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT58), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n834), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n732), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n835), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n851), .B1(new_n858), .B2(new_n850), .ZN(G1344gat));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n432), .A3(new_n316), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n809), .A2(new_n810), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n847), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n846), .A2(new_n684), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(KEYINPUT57), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n865), .A2(new_n316), .A3(new_n731), .A4(new_n834), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n432), .C1(new_n849), .C2(new_n316), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n860), .B1(new_n867), .B2(new_n868), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n855), .A2(new_n437), .A3(new_n242), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n849), .A2(new_n242), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n437), .B2(new_n871), .ZN(G1346gat));
  AND2_X1   g671(.A1(new_n849), .A2(new_n295), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n822), .A2(new_n438), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n873), .A2(new_n438), .B1(new_n854), .B2(new_n874), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n674), .A2(new_n629), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n862), .A2(new_n632), .A3(new_n595), .A4(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(G169gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(new_n878), .A3(new_n669), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n732), .A2(new_n588), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT121), .B1(new_n811), .B2(new_n629), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n862), .A2(new_n882), .A3(new_n517), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n345), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n879), .B1(new_n885), .B2(new_n878), .ZN(G1348gat));
  OAI21_X1  g685(.A(G176gat), .B1(new_n877), .B2(new_n689), .ZN(new_n887));
  INV_X1    g686(.A(new_n884), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n689), .A2(G176gat), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(G1349gat));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n242), .A2(new_n391), .A3(new_n393), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G183gat), .B1(new_n877), .B2(new_n243), .ZN(new_n894));
  AND2_X1   g693(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n891), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n897), .B2(KEYINPUT122), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n891), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n877), .B2(new_n688), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT61), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n384), .A3(new_n295), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1351gat));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n846), .B2(new_n684), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n862), .A2(new_n847), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n876), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n680), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n345), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G197gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n680), .A2(new_n731), .A3(new_n632), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n881), .B2(new_n883), .ZN(new_n916));
  INV_X1    g715(.A(G197gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n345), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(new_n316), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n316), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G204gat), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n925), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n348), .A3(new_n242), .ZN(new_n932));
  OR2_X1    g731(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n242), .B(new_n909), .C1(new_n905), .C2(new_n906), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n348), .B1(new_n935), .B2(KEYINPUT126), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n865), .A2(KEYINPUT126), .A3(new_n242), .A4(new_n909), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n940), .A2(new_n938), .A3(G211gat), .A4(new_n933), .ZN(new_n941));
  NAND2_X1  g740(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n932), .B1(new_n939), .B2(new_n943), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n916), .B2(new_n295), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n688), .A2(new_n356), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n911), .B2(new_n946), .ZN(G1355gat));
endmodule


