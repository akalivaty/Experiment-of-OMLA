//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1037, new_n1038;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT23), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n210), .A2(KEYINPUT23), .A3(new_n204), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(G183gat), .B(G190gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT25), .B(new_n220), .C1(new_n222), .C2(new_n207), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n226), .B1(new_n231), .B2(KEYINPUT24), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n220), .A2(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n232), .A2(KEYINPUT65), .A3(new_n209), .A4(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n224), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(KEYINPUT27), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT27), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n239), .A3(new_n229), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n207), .A2(KEYINPUT26), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n204), .A2(new_n205), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT26), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G169gat), .B2(G176gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n243), .B(new_n225), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n241), .ZN(new_n249));
  INV_X1    g048(.A(new_n236), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G113gat), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G120gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G127gat), .B(G134gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G127gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G134gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n265), .C1(new_n266), .C2(KEYINPUT1), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n254), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n264), .A2(KEYINPUT1), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n259), .A2(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n267), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n271), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n235), .A2(new_n251), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT33), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G15gat), .B(G43gat), .Z(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n286), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n280), .B(KEYINPUT32), .C1(new_n282), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n275), .B1(new_n274), .B2(new_n279), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n287), .B2(new_n289), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n290), .A2(new_n291), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n296));
  NOR3_X1   g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n289), .ZN(new_n299));
  INV_X1    g098(.A(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n287), .A2(new_n289), .A3(new_n292), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n202), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n296), .B1(new_n293), .B2(new_n294), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n302), .A3(new_n298), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT36), .ZN(new_n307));
  XOR2_X1   g106(.A(G1gat), .B(G29gat), .Z(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT74), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(G141gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(G148gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G155gat), .ZN(new_n325));
  INV_X1    g124(.A(G155gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n313), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(G148gat), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n332), .B2(new_n319), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n336), .B2(new_n324), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n323), .A2(new_n328), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n273), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n273), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT5), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(new_n273), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n345), .B1(new_n338), .B2(new_n273), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n278), .B1(new_n338), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n322), .A2(new_n318), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n321), .B1(new_n319), .B2(new_n320), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n328), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n337), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n343), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT77), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n343), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n355), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n273), .B1(new_n361), .B2(KEYINPUT3), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n339), .A2(KEYINPUT4), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n346), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n344), .B1(new_n359), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(KEYINPUT3), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n278), .A3(new_n356), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n339), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n370), .B(new_n371), .C1(new_n365), .C2(KEYINPUT79), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n360), .A2(KEYINPUT5), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n312), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT5), .ZN(new_n377));
  INV_X1    g176(.A(new_n341), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n339), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n379), .B2(new_n360), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n366), .B1(new_n363), .B2(new_n365), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n312), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n347), .A2(KEYINPUT79), .A3(new_n348), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n371), .ZN(new_n386));
  OR3_X1    g185(.A1(new_n385), .A2(new_n386), .A3(new_n374), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT6), .B(new_n312), .C1(new_n368), .C2(new_n375), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G8gat), .B(G36gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT73), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n249), .A2(new_n250), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n398), .A2(new_n247), .A3(new_n242), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n229), .A2(G183gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n227), .A2(G190gat), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT24), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n233), .A2(new_n402), .A3(new_n215), .A4(new_n209), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n209), .A3(new_n212), .A4(new_n215), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n219), .A2(new_n403), .B1(new_n404), .B2(new_n203), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n405), .B2(new_n234), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n397), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  AND2_X1   g206(.A1(G211gat), .A2(G218gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(G211gat), .A2(G218gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(G197gat), .A2(G204gat), .ZN(new_n411));
  NOR2_X1   g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G211gat), .B(G218gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G197gat), .B(G204gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n414), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT71), .B(new_n410), .C1(new_n413), .C2(new_n414), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n397), .B1(new_n235), .B2(new_n251), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n397), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n252), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n406), .B2(new_n397), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(KEYINPUT72), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n396), .B(new_n427), .C1(new_n434), .C2(new_n424), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n427), .B1(new_n434), .B2(new_n424), .ZN(new_n438));
  INV_X1    g237(.A(new_n396), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT72), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n431), .B(new_n397), .C1(new_n235), .C2(new_n251), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n407), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n423), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(KEYINPUT30), .A3(new_n396), .A4(new_n427), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n392), .A2(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT80), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n421), .A2(new_n429), .A3(new_n422), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT81), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n421), .A2(new_n456), .A3(new_n429), .A4(new_n422), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n350), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n361), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT82), .ZN(new_n460));
  NAND2_X1  g259(.A1(G228gat), .A2(G233gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n356), .A2(new_n429), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n424), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT29), .B1(new_n338), .B2(new_n350), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT83), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(new_n468), .A3(new_n361), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G22gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n424), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n415), .A2(new_n419), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT3), .B1(new_n473), .B2(new_n429), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(new_n338), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n461), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n471), .B1(new_n470), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n453), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G22gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n470), .A2(new_n471), .A3(new_n476), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n452), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n304), .A2(new_n307), .B1(new_n448), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n360), .C1(new_n385), .C2(new_n386), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n384), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT39), .B1(new_n379), .B2(new_n360), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n372), .B2(new_n360), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n360), .B1(new_n385), .B2(new_n386), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n488), .B1(new_n342), .B2(new_n343), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(KEYINPUT40), .A3(new_n384), .A4(new_n489), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n493), .A2(new_n376), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n498), .A2(new_n446), .B1(new_n483), .B2(new_n479), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n430), .A2(new_n423), .A3(new_n425), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n423), .B2(new_n443), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT37), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n396), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n443), .A2(new_n424), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n430), .A2(new_n425), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(new_n423), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT38), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n503), .A2(new_n507), .B1(new_n396), .B2(new_n501), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n439), .B1(new_n438), .B2(KEYINPUT37), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n501), .A2(new_n502), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n508), .A2(new_n511), .A3(new_n391), .A4(new_n390), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n484), .A2(new_n305), .A3(new_n306), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT35), .B1(new_n514), .B2(new_n448), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n305), .A2(new_n306), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n446), .B1(new_n391), .B2(new_n390), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n484), .A4(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n486), .A2(new_n513), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  INV_X1    g324(.A(G1gat), .ZN(new_n526));
  INV_X1    g325(.A(G15gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(G22gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n471), .A2(G15gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n531), .B(G8gat), .C1(new_n525), .C2(new_n524), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n522), .B(new_n536), .C1(new_n523), .C2(G1gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT14), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G43gat), .ZN(new_n549));
  INV_X1    g348(.A(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n552));
  NAND2_X1  g351(.A1(G43gat), .A2(G50gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n541), .A2(new_n548), .A3(KEYINPUT15), .A4(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n554), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(KEYINPUT15), .B2(new_n540), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n541), .A2(KEYINPUT15), .A3(new_n554), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n562), .B(new_n557), .C1(KEYINPUT15), .C2(new_n540), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n532), .A2(new_n538), .A3(new_n563), .A4(new_n555), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT13), .Z(new_n567));
  INV_X1    g366(.A(new_n539), .ZN(new_n568));
  INV_X1    g367(.A(new_n559), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(KEYINPUT89), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(KEYINPUT86), .A2(KEYINPUT17), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT86), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n563), .A2(new_n573), .A3(new_n574), .A4(new_n555), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n539), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n566), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n532), .A2(new_n538), .B1(new_n563), .B2(new_n555), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n571), .B1(new_n581), .B2(KEYINPUT18), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT18), .ZN(new_n583));
  NOR4_X1   g382(.A1(new_n578), .A2(new_n583), .A3(new_n579), .A4(new_n580), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n521), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G113gat), .B(G141gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(G197gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT11), .B(G169gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT12), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n521), .B(new_n590), .C1(new_n582), .C2(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR3_X1   g393(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT90), .B1(G71gat), .B2(G78gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  AOI211_X1 g398(.A(new_n595), .B(new_n598), .C1(new_n599), .C2(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G57gat), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n601), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n602));
  OAI21_X1  g401(.A(G64gat), .B1(new_n601), .B2(KEYINPUT91), .ZN(new_n603));
  INV_X1    g402(.A(G71gat), .ZN(new_n604));
  INV_X1    g403(.A(G78gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT9), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n602), .A2(new_n603), .B1(new_n597), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n262), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n568), .B1(new_n610), .B2(new_n609), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G155gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n616), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(G85gat), .B2(G92gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT92), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(KEYINPUT7), .A3(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT8), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n630), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT93), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n628), .B(new_n632), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G99gat), .B(G106gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n622), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n631), .A2(KEYINPUT7), .A3(new_n625), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT7), .B1(new_n631), .B2(new_n625), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(new_n645), .A3(KEYINPUT94), .A4(new_n639), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n638), .A2(new_n640), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n638), .A2(KEYINPUT95), .A3(new_n640), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n576), .A2(new_n577), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n569), .ZN(new_n657));
  AND3_X1   g456(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G190gat), .B(G218gat), .Z(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n654), .A2(new_n655), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT96), .B1(new_n652), .B2(new_n653), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n659), .B(new_n666), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n662), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n665), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(new_n656), .B2(new_n659), .ZN(new_n672));
  INV_X1    g471(.A(new_n669), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n642), .A2(new_n645), .A3(new_n639), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n648), .A2(new_n678), .A3(new_n608), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT97), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n678), .A2(new_n648), .A3(new_n608), .A4(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n652), .A2(new_n609), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n677), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT98), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n685), .A2(new_n687), .B1(new_n686), .B2(new_n683), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n652), .A2(new_n609), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n680), .A2(new_n682), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n684), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n677), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n686), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n686), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n692), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n688), .A2(new_n692), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n621), .A2(new_n675), .A3(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n520), .A2(new_n594), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n392), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT99), .B(G1gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1324gat));
  XOR2_X1   g506(.A(KEYINPUT16), .B(G8gat), .Z(new_n708));
  AND3_X1   g507(.A1(new_n703), .A2(new_n446), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n533), .B1(new_n703), .B2(new_n446), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT42), .B2(new_n709), .ZN(G1325gat));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n527), .A3(new_n516), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n304), .A2(new_n307), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(new_n527), .ZN(G1326gat));
  NAND2_X1  g516(.A1(new_n703), .A2(new_n485), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT100), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  NAND2_X1  g520(.A1(new_n515), .A2(new_n519), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n448), .A2(new_n485), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n714), .A2(new_n513), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n675), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n698), .A2(new_n700), .ZN(new_n726));
  INV_X1    g525(.A(new_n687), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n699), .B1(new_n697), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n728), .B2(new_n691), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n621), .A2(new_n594), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n542), .A3(new_n704), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT101), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT44), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n520), .B2(new_n675), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n724), .ZN(new_n738));
  INV_X1    g537(.A(new_n675), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n737), .A2(new_n741), .A3(new_n730), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n704), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n734), .B1(new_n542), .B2(new_n743), .ZN(G1328gat));
  NAND3_X1  g543(.A1(new_n731), .A2(new_n543), .A3(new_n446), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT46), .Z(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n446), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G36gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(G1329gat));
  NAND3_X1  g550(.A1(new_n742), .A2(G43gat), .A3(new_n715), .ZN(new_n752));
  INV_X1    g551(.A(new_n731), .ZN(new_n753));
  INV_X1    g552(.A(new_n516), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n549), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g556(.A1(new_n742), .A2(G50gat), .A3(new_n485), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n550), .B1(new_n753), .B2(new_n484), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g560(.A(new_n621), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n594), .A2(new_n729), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n520), .A2(new_n762), .A3(new_n739), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n704), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n446), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  AOI21_X1  g569(.A(new_n604), .B1(new_n764), .B2(new_n715), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n754), .A2(G71gat), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n764), .A2(new_n485), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  OAI21_X1  g575(.A(KEYINPUT105), .B1(new_n520), .B2(new_n675), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n738), .A2(new_n778), .A3(new_n739), .ZN(new_n779));
  INV_X1    g578(.A(new_n594), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n621), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n781), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n725), .B2(new_n778), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(KEYINPUT51), .A3(new_n777), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(new_n629), .A3(new_n704), .A4(new_n729), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n621), .A2(new_n763), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n737), .A2(new_n741), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT104), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n737), .A2(new_n741), .A3(new_n793), .A4(new_n790), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n704), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n789), .B1(new_n629), .B2(new_n795), .ZN(G1336gat));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n737), .A2(new_n741), .A3(new_n446), .A4(new_n790), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n798), .B2(G92gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n447), .A2(new_n701), .A3(G92gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n784), .B2(new_n787), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n799), .B1(new_n802), .B2(KEYINPUT107), .ZN(new_n803));
  AND4_X1   g602(.A1(KEYINPUT51), .A2(new_n777), .A3(new_n779), .A4(new_n781), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n786), .B2(new_n777), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n446), .A3(new_n794), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n782), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n783), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n782), .A2(new_n813), .A3(KEYINPUT51), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n800), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n810), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n797), .B1(new_n809), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n807), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n802), .A2(KEYINPUT107), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n799), .ZN(new_n822));
  AOI211_X1 g621(.A(KEYINPUT106), .B(new_n783), .C1(new_n786), .C2(new_n777), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT51), .B1(new_n782), .B2(new_n813), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n825), .A2(new_n800), .B1(new_n811), .B2(G92gat), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(KEYINPUT108), .C1(new_n826), .C2(new_n810), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n827), .ZN(G1337gat));
  NAND3_X1  g627(.A1(new_n792), .A2(new_n715), .A3(new_n794), .ZN(new_n829));
  XOR2_X1   g628(.A(KEYINPUT109), .B(G99gat), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n754), .A2(new_n701), .A3(new_n830), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT110), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n788), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(G1338gat));
  NOR3_X1   g634(.A1(new_n484), .A2(G106gat), .A3(new_n701), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n815), .A2(new_n816), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n825), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n792), .A2(new_n485), .A3(new_n794), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G106gat), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n791), .A2(new_n484), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n845), .B2(G106gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n788), .A2(new_n836), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(G1339gat));
  NOR2_X1   g648(.A1(new_n702), .A2(new_n780), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n685), .A2(new_n687), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n691), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n686), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n685), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n697), .A2(new_n727), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n852), .B1(new_n697), .B2(new_n686), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n685), .A2(new_n687), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT112), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n582), .A2(new_n584), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n565), .A2(new_n570), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n580), .B1(new_n653), .B2(new_n568), .ZN(new_n867));
  OAI22_X1  g666(.A1(new_n866), .A2(new_n567), .B1(new_n566), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n865), .A2(new_n590), .B1(new_n589), .B2(new_n868), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n670), .A2(new_n674), .A3(new_n726), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n857), .B1(new_n855), .B2(new_n856), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n859), .A2(KEYINPUT112), .A3(new_n860), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n863), .B(new_n691), .C1(new_n851), .C2(new_n852), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n864), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n867), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n583), .B1(new_n877), .B2(new_n579), .ZN(new_n878));
  INV_X1    g677(.A(new_n584), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n878), .A2(new_n590), .A3(new_n879), .A4(new_n571), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n868), .A2(new_n589), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT113), .B1(new_n701), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n729), .A2(new_n884), .A3(new_n869), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n592), .A2(new_n593), .A3(new_n726), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n873), .B2(new_n874), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n864), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n876), .B1(new_n889), .B2(new_n739), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n850), .B1(new_n890), .B2(new_n762), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n514), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n392), .A2(new_n446), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n780), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n729), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g697(.A1(new_n894), .A2(new_n621), .ZN(new_n899));
  NOR2_X1   g698(.A1(KEYINPUT114), .A2(G127gat), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n899), .B(new_n900), .Z(G1342gat));
  AND3_X1   g700(.A1(new_n892), .A2(new_n739), .A3(new_n893), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n260), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT56), .Z(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n260), .B2(new_n902), .ZN(G1343gat));
  INV_X1    g704(.A(new_n850), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n864), .A2(new_n870), .A3(new_n875), .ZN(new_n907));
  INV_X1    g706(.A(new_n887), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n875), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT55), .B1(new_n873), .B2(new_n853), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n883), .B(new_n885), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n911), .B2(new_n675), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n912), .B2(new_n621), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n485), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n714), .A2(new_n893), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n914), .A2(G141gat), .A3(new_n594), .A4(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n891), .B2(new_n484), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n864), .A2(new_n888), .B1(new_n729), .B2(new_n869), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n876), .B1(new_n919), .B2(new_n739), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n850), .B1(new_n920), .B2(new_n762), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n484), .A2(new_n917), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT115), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n909), .A2(new_n910), .B1(new_n701), .B2(new_n882), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n675), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n621), .B1(new_n927), .B2(new_n876), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n925), .B(new_n922), .C1(new_n928), .C2(new_n850), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n915), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n780), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n330), .A2(new_n331), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n916), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n935));
  NOR2_X1   g734(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n936));
  AND2_X1   g735(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(G1344gat));
  NAND3_X1  g738(.A1(new_n913), .A2(KEYINPUT117), .A3(new_n922), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n891), .B2(new_n923), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n917), .B1(new_n921), .B2(new_n484), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n729), .A3(new_n931), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n913), .A2(new_n485), .A3(new_n931), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT59), .B1(new_n947), .B2(new_n701), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n701), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n315), .A2(new_n948), .B1(new_n930), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT118), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n946), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1345gat));
  NAND2_X1  g754(.A1(new_n930), .A2(new_n931), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(new_n762), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n621), .A2(new_n336), .ZN(new_n958));
  OAI22_X1  g757(.A1(new_n957), .A2(new_n336), .B1(new_n947), .B2(new_n958), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n956), .B2(new_n675), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n675), .A2(G162gat), .A3(new_n446), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n714), .A2(new_n961), .A3(new_n704), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n914), .B2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n704), .A2(new_n447), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n891), .A2(new_n514), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n780), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT119), .A3(G169gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT119), .B1(new_n967), .B2(G169gat), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n968), .A2(new_n969), .B1(G169gat), .B2(new_n967), .ZN(G1348gat));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n971));
  AOI21_X1  g770(.A(G176gat), .B1(new_n966), .B2(new_n729), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n210), .A2(new_n211), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n966), .A2(new_n975), .A3(new_n729), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n976), .A2(KEYINPUT121), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(KEYINPUT121), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n971), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n974), .A2(new_n977), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n983), .A2(KEYINPUT122), .A3(new_n979), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1349gat));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n986));
  INV_X1    g785(.A(new_n514), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n913), .A2(new_n987), .A3(new_n621), .A4(new_n964), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n227), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n237), .A2(new_n239), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n986), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT124), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n892), .A2(new_n991), .A3(new_n621), .A4(new_n964), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n989), .A2(new_n996), .A3(KEYINPUT123), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT60), .A4(new_n997), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n989), .A2(new_n996), .A3(KEYINPUT123), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT123), .B1(new_n989), .B2(new_n996), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT60), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n990), .B2(new_n993), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT124), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n998), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(new_n1005), .ZN(G1350gat));
  NOR2_X1   g805(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n966), .B2(new_n739), .ZN(new_n1008));
  NAND2_X1  g807(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1008), .B(new_n1009), .Z(G1351gat));
  XOR2_X1   g809(.A(KEYINPUT125), .B(G197gat), .Z(new_n1011));
  NOR2_X1   g810(.A1(new_n715), .A2(new_n965), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n944), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1011), .B1(new_n1013), .B2(new_n594), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n714), .A2(new_n485), .A3(new_n964), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n891), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n594), .A2(new_n1011), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(G1352gat));
  OAI21_X1  g818(.A(G204gat), .B1(new_n1013), .B2(new_n701), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n701), .A2(G204gat), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g821(.A(new_n1022), .B(KEYINPUT62), .Z(new_n1023));
  NAND2_X1  g822(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1024), .A2(KEYINPUT126), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1025), .A2(new_n1027), .ZN(G1353gat));
  OR3_X1    g827(.A1(new_n1017), .A2(G211gat), .A3(new_n762), .ZN(new_n1029));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n944), .A2(new_n621), .A3(new_n1012), .ZN(new_n1031));
  AND4_X1   g830(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1032));
  OAI21_X1  g831(.A(G211gat), .B1(new_n1030), .B2(KEYINPUT63), .ZN(new_n1033));
  INV_X1    g832(.A(new_n1033), .ZN(new_n1034));
  AOI22_X1  g833(.A1(new_n1031), .A2(new_n1034), .B1(new_n1030), .B2(KEYINPUT63), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1029), .B1(new_n1032), .B2(new_n1035), .ZN(G1354gat));
  OAI21_X1  g835(.A(G218gat), .B1(new_n1013), .B2(new_n675), .ZN(new_n1037));
  OR3_X1    g836(.A1(new_n1017), .A2(G218gat), .A3(new_n675), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1037), .A2(new_n1038), .ZN(G1355gat));
endmodule


