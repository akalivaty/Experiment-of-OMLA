//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT30), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n211), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT67), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT27), .B(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT28), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n215), .A2(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n211), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT64), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n224), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n240), .A2(new_n241), .B1(new_n226), .B2(new_n225), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n243), .A3(KEYINPUT66), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n227), .A2(new_n228), .B1(new_n207), .B2(new_n230), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n211), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n238), .A2(new_n242), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n223), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G226gat), .A2(G233gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n215), .A2(new_n216), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n221), .A2(new_n222), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n252), .B2(new_n253), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n255), .A2(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  INV_X1    g063(.A(G211gat), .ZN(new_n265));
  INV_X1    g064(.A(G218gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n264), .B1(KEYINPUT22), .B2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n256), .B1(new_n255), .B2(KEYINPUT29), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n275), .B(new_n256), .C1(new_n255), .C2(KEYINPUT29), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n257), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n272), .B1(new_n278), .B2(new_n271), .ZN(new_n279));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  NOR2_X1   g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n284), .B(new_n272), .C1(new_n278), .C2(new_n271), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n204), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G120gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT68), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n287), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g098(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(G120gat), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n299), .B1(new_n289), .B2(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(new_n297), .A2(new_n303), .A3(KEYINPUT70), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT70), .ZN(new_n305));
  INV_X1    g104(.A(new_n287), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n298), .B1(new_n295), .B2(KEYINPUT68), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n293), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n289), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n298), .A3(new_n287), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n305), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G148gat), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(G141gat), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G155gat), .ZN(new_n321));
  INV_X1    g120(.A(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n323), .A2(new_n325), .ZN(new_n330));
  INV_X1    g129(.A(G141gat), .ZN(new_n331));
  INV_X1    g130(.A(G148gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n326), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n314), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n316), .A2(new_n319), .B1(new_n324), .B2(new_n327), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  NOR3_X1   g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT77), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT4), .B1(new_n313), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n297), .B2(new_n303), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n309), .A2(KEYINPUT76), .A3(new_n311), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n346), .A3(new_n336), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(new_n338), .B2(new_n339), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT4), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n297), .A2(new_n303), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n338), .A2(new_n339), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n349), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n342), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(KEYINPUT5), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n349), .A2(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n313), .A2(new_n341), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n352), .A2(new_n350), .A3(new_n309), .A4(new_n311), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT78), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n351), .A2(new_n365), .A3(new_n350), .A4(new_n352), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n360), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  INV_X1    g168(.A(new_n352), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n344), .A3(new_n345), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n353), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n357), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n359), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G1gat), .B(G29gat), .Z(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G57gat), .B(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n375), .B2(new_n380), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n350), .B1(new_n313), .B2(new_n341), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n364), .A2(new_n366), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n356), .B(new_n349), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n386), .A2(new_n373), .B1(new_n355), .B2(new_n358), .ZN(new_n387));
  INV_X1    g186(.A(new_n380), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n381), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n204), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n279), .A2(new_n282), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n391), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n286), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT81), .Z(new_n398));
  XNOR2_X1  g197(.A(new_n268), .B(new_n269), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n341), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n352), .B2(new_n346), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(new_n399), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n398), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT82), .B(G22gat), .ZN(new_n406));
  OAI211_X1 g205(.A(G228gat), .B(G233gat), .C1(new_n401), .C2(new_n352), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n405), .B(new_n406), .C1(new_n404), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n398), .ZN(new_n409));
  OR2_X1    g208(.A1(new_n403), .A2(new_n399), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n346), .B1(new_n271), .B2(KEYINPUT29), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n337), .B2(new_n340), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n407), .A2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(G22gat), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT31), .B(G50gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n408), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n418), .B(KEYINPUT80), .Z(new_n421));
  INV_X1    g220(.A(new_n406), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n413), .B2(new_n414), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n408), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n396), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT36), .ZN(new_n427));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT66), .B1(new_n236), .B2(new_n243), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n252), .A2(new_n253), .A3(new_n245), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n260), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n312), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n309), .A2(new_n305), .A3(new_n311), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n255), .A2(new_n313), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n430), .B1(new_n440), .B2(KEYINPUT33), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT32), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n439), .ZN(new_n445));
  INV_X1    g244(.A(new_n431), .ZN(new_n446));
  AOI221_X4 g245(.A(new_n442), .B1(KEYINPUT33), .B2(new_n430), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT71), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n438), .A2(new_n439), .A3(new_n431), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT34), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n444), .A2(new_n451), .A3(new_n447), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n449), .B(KEYINPUT34), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n434), .A2(new_n437), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n255), .A2(new_n313), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT32), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n459), .A3(new_n430), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n443), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n453), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n448), .B1(new_n452), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n453), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n427), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n451), .B1(new_n444), .B2(new_n447), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n461), .A3(new_n453), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n426), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT86), .B1(new_n387), .B2(new_n388), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n375), .A2(new_n473), .A3(new_n380), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n355), .A2(new_n356), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT84), .B(KEYINPUT39), .Z(new_n478));
  AOI21_X1  g277(.A(new_n380), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n371), .A2(new_n353), .A3(new_n356), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT85), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(KEYINPUT39), .C1(new_n356), .C2(new_n355), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g282(.A1(new_n479), .A2(new_n476), .A3(new_n482), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n475), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n273), .A2(KEYINPUT72), .B1(new_n257), .B2(new_n261), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n399), .B1(new_n486), .B2(new_n276), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n284), .B1(new_n487), .B2(new_n272), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n391), .B1(new_n392), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n204), .B1(new_n285), .B2(new_n393), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT83), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n286), .A2(new_n492), .A3(new_n395), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n485), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT6), .B1(new_n387), .B2(new_n388), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n496), .A3(new_n474), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n381), .A3(new_n392), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n274), .A2(new_n399), .A3(new_n276), .A4(new_n277), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n261), .A2(new_n262), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n271), .C1(new_n434), .C2(new_n256), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n505), .A3(new_n399), .A4(new_n276), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT37), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n282), .A2(KEYINPUT38), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n279), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n498), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n284), .B1(new_n279), .B2(new_n511), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(KEYINPUT89), .B(new_n284), .C1(new_n279), .C2(new_n511), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n279), .A2(new_n511), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT38), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n425), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n471), .B1(new_n495), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n425), .B1(new_n463), .B2(new_n465), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n286), .A2(new_n390), .A3(new_n395), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n525), .B1(new_n420), .B2(new_n424), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n497), .B2(new_n381), .ZN(new_n530));
  AND4_X1   g329(.A1(new_n491), .A2(new_n493), .A3(new_n530), .A4(new_n469), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n202), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n467), .A2(new_n468), .B1(KEYINPUT71), .B2(new_n464), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n464), .A2(KEYINPUT71), .A3(new_n453), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT36), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n469), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n427), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n536), .A2(new_n538), .B1(new_n425), .B2(new_n396), .ZN(new_n539));
  INV_X1    g338(.A(new_n425), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT38), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n519), .A2(new_n520), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n517), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n508), .A2(new_n512), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(new_n381), .A3(new_n392), .A4(new_n497), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n540), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n539), .B1(new_n546), .B2(new_n494), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n547), .B(KEYINPUT90), .C1(new_n528), .C2(new_n531), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT91), .B(G29gat), .Z(new_n550));
  XOR2_X1   g349(.A(KEYINPUT92), .B(G36gat), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g353(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(KEYINPUT15), .A3(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n555), .A2(new_n562), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n554), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n558), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT17), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  AND2_X1   g367(.A1(KEYINPUT94), .A2(G1gat), .ZN(new_n569));
  OAI21_X1  g368(.A(KEYINPUT16), .B1(KEYINPUT94), .B2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(KEYINPUT95), .C1(G1gat), .C2(new_n568), .ZN(new_n572));
  INV_X1    g371(.A(G8gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n566), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT18), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n576), .A4(new_n578), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n574), .B(new_n566), .Z(new_n583));
  XOR2_X1   g382(.A(new_n576), .B(KEYINPUT13), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G197gat), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT11), .B(G169gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT12), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n581), .A2(new_n593), .A3(new_n582), .A4(new_n585), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n592), .A2(KEYINPUT96), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT96), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  OAI211_X1 g398(.A(G85gat), .B(G92gat), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(KEYINPUT99), .B2(KEYINPUT7), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n600), .B(KEYINPUT100), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(new_n598), .A3(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT8), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(G85gat), .B2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT101), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n603), .A2(new_n605), .A3(new_n613), .A4(new_n609), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n566), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT41), .ZN(new_n616));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n614), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n567), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n616), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(G71gat), .A2(G78gat), .ZN(new_n631));
  NOR2_X1   g430(.A1(G71gat), .A2(G78gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G57gat), .B(G64gat), .Z(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(KEYINPUT97), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(KEYINPUT9), .B2(new_n631), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(G127gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n577), .B1(KEYINPUT21), .B2(new_n639), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G155gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n630), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT102), .ZN(new_n656));
  INV_X1    g455(.A(new_n639), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n619), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n612), .A2(new_n639), .A3(new_n614), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n660), .A2(new_n659), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n658), .A2(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n665), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n661), .A2(new_n662), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n664), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n670), .ZN(new_n677));
  INV_X1    g476(.A(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n655), .A2(new_n656), .A3(new_n681), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n549), .A2(new_n597), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n390), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(G1gat), .Z(G1324gat));
  INV_X1    g484(.A(new_n493), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n492), .B1(new_n286), .B2(new_n395), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G8gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n573), .B2(new_n689), .ZN(new_n693));
  MUX2_X1   g492(.A(new_n692), .B(new_n693), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g493(.A1(new_n466), .A2(new_n470), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n683), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n537), .A2(G15gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n683), .B2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n540), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT105), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n549), .A2(new_n597), .ZN(new_n704));
  INV_X1    g503(.A(new_n653), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n629), .A4(new_n681), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(new_n390), .A3(new_n550), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT45), .Z(new_n708));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n528), .B2(new_n531), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n540), .B1(new_n534), .B2(new_n535), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT35), .B1(new_n711), .B2(new_n396), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n491), .A2(new_n493), .A3(new_n530), .A4(new_n469), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n547), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n629), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n630), .A2(new_n717), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n533), .A2(new_n548), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n680), .B(KEYINPUT107), .Z(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n592), .A2(new_n594), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n722), .A2(new_n653), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n550), .B1(new_n727), .B2(new_n390), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n728), .ZN(G1328gat));
  NOR3_X1   g528(.A1(new_n706), .A2(new_n688), .A3(new_n551), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT46), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n551), .B1(new_n727), .B2(new_n688), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1329gat));
  NOR2_X1   g532(.A1(new_n706), .A2(new_n537), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n695), .A2(G43gat), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n734), .A2(G43gat), .B1(new_n727), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g536(.A(G50gat), .B1(new_n727), .B2(new_n540), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n738), .B2(KEYINPUT109), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n540), .A2(G50gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n706), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n739), .B(new_n741), .ZN(G1331gat));
  AND4_X1   g541(.A1(new_n656), .A2(new_n655), .A3(new_n722), .A4(new_n725), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n715), .ZN(new_n744));
  INV_X1    g543(.A(new_n390), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  INV_X1    g546(.A(new_n688), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT49), .B(G64gat), .Z(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(G1333gat));
  NAND3_X1  g551(.A1(new_n744), .A2(G71gat), .A3(new_n695), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT110), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n744), .A2(new_n469), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(G71gat), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n744), .A2(new_n425), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  XNOR2_X1  g558(.A(new_n723), .B(KEYINPUT106), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n653), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n680), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT111), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n718), .A2(new_n720), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n390), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n715), .A2(new_n629), .A3(new_n761), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n715), .A2(KEYINPUT51), .A3(new_n629), .A4(new_n761), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n681), .A2(G85gat), .A3(new_n390), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT112), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n766), .B1(new_n772), .B2(new_n774), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n688), .A2(G92gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n771), .A2(new_n722), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n718), .A2(new_n748), .A3(new_n720), .A4(new_n763), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n721), .B1(new_n769), .B2(new_n770), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n786), .A2(new_n777), .B1(new_n779), .B2(G92gat), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n787), .B2(new_n781), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT113), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n776), .B(new_n785), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n784), .B1(new_n787), .B2(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n782), .A2(new_n783), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n776), .B1(new_n795), .B2(new_n785), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n792), .A2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n765), .B2(new_n696), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n681), .A2(G99gat), .A3(new_n537), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n772), .B2(new_n799), .ZN(G1338gat));
  NAND2_X1  g599(.A1(new_n764), .A2(new_n425), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n803), .A3(new_n425), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n802), .B2(KEYINPUT116), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n808), .A3(new_n804), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n807), .B1(new_n806), .B2(new_n809), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(G1339gat));
  AOI21_X1  g611(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n583), .A2(new_n584), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n590), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n594), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n680), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n678), .B1(new_n676), .B2(KEYINPUT54), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n666), .A2(new_n667), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT54), .B1(new_n675), .B2(new_n664), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n819), .B(KEYINPUT55), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n674), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n817), .B1(new_n826), .B2(new_n725), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT118), .B(new_n817), .C1(new_n826), .C2(new_n725), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n630), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n826), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n629), .A3(new_n816), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n653), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n682), .A2(new_n760), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n540), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n748), .A2(new_n537), .ZN(new_n838));
  INV_X1    g637(.A(new_n597), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(new_n745), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT119), .B1(new_n840), .B2(G113gat), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n534), .A2(new_n535), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n748), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n837), .A2(new_n745), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n760), .A2(new_n300), .A3(new_n301), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n842), .A2(new_n843), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n288), .A3(new_n680), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n837), .A2(new_n745), .A3(new_n838), .A4(new_n722), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(KEYINPUT120), .A3(G120gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT120), .B1(new_n851), .B2(G120gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n846), .A2(new_n643), .A3(new_n653), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n745), .A3(new_n838), .ZN(new_n857));
  OAI21_X1  g656(.A(G127gat), .B1(new_n857), .B2(new_n705), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1342gat));
  XOR2_X1   g658(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n630), .A2(G134gat), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n847), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n857), .B2(new_n630), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n862), .A3(new_n860), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  INV_X1    g667(.A(new_n315), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n425), .C1(new_n834), .C2(new_n835), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n748), .A2(new_n390), .A3(new_n695), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n825), .A2(new_n674), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n597), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT55), .B1(new_n822), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n819), .B(KEYINPUT122), .C1(new_n820), .C2(new_n821), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT123), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n821), .B1(new_n666), .B2(new_n667), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(new_n818), .ZN(new_n880));
  AND4_X1   g679(.A1(KEYINPUT123), .A2(new_n877), .A3(new_n880), .A4(new_n823), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n874), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n629), .B1(new_n882), .B2(new_n817), .ZN(new_n883));
  INV_X1    g682(.A(new_n833), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n705), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n835), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n540), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n871), .B(new_n872), .C1(new_n887), .C2(new_n870), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n869), .B1(new_n888), .B2(new_n725), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n597), .A2(G141gat), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n836), .A2(new_n425), .A3(new_n872), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n868), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n868), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n885), .A2(new_n886), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n540), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n895), .A2(new_n839), .A3(new_n871), .A4(new_n872), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n896), .B2(new_n869), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n893), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n869), .B1(new_n888), .B2(new_n597), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  INV_X1    g701(.A(new_n891), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n895), .A2(new_n760), .A3(new_n871), .A4(new_n872), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n869), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n901), .B(new_n902), .C1(new_n905), .C2(new_n868), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n898), .A2(new_n906), .ZN(G1344gat));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n836), .A2(new_n425), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n832), .A2(new_n629), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT125), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n816), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n883), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n653), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n682), .A2(new_n839), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n870), .B(new_n425), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n910), .A2(new_n680), .A3(new_n872), .A4(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n908), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n888), .A2(new_n681), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n317), .A2(new_n318), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n836), .A2(new_n425), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n872), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n680), .A2(new_n923), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n920), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n888), .B2(new_n705), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n653), .A2(new_n321), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(G1346gat));
  OAI21_X1  g730(.A(G162gat), .B1(new_n888), .B2(new_n630), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n629), .A2(new_n322), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n926), .B2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n688), .A2(new_n745), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n537), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n837), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n205), .A3(new_n597), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n836), .A2(new_n526), .A3(new_n935), .ZN(new_n940));
  AOI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n760), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n939), .A2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n938), .B2(new_n721), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n206), .A3(new_n680), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n938), .B2(new_n705), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n217), .A3(new_n653), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n940), .A2(new_n218), .A3(new_n629), .ZN(new_n953));
  OAI21_X1  g752(.A(G190gat), .B1(new_n938), .B2(new_n630), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  AND2_X1   g756(.A1(new_n910), .A2(new_n918), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n936), .A2(new_n695), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(G197gat), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n597), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n925), .A2(new_n959), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n925), .A2(KEYINPUT126), .A3(new_n959), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n760), .A3(new_n967), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n961), .A2(new_n963), .B1(new_n968), .B2(new_n962), .ZN(G1352gat));
  OAI21_X1  g768(.A(G204gat), .B1(new_n960), .B2(new_n721), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n681), .A2(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n925), .A2(new_n959), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT62), .Z(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(new_n973), .ZN(G1353gat));
  NAND4_X1  g773(.A1(new_n910), .A2(new_n653), .A3(new_n918), .A4(new_n959), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n966), .A2(new_n967), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n653), .A2(new_n265), .ZN(new_n979));
  OAI22_X1  g778(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n960), .B2(new_n630), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n266), .A3(new_n629), .A4(new_n967), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


