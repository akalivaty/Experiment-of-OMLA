//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G116), .ZN(new_n214));
  INV_X1    g0014(.A(G270), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT65), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n216), .A2(new_n217), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G97), .A2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n207), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n226), .B1(KEYINPUT66), .B2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n203), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n210), .B(new_n229), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n215), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n212), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n230), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n231), .A2(KEYINPUT68), .A3(G33), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n202), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n262), .A2(new_n212), .B1(new_n231), .B2(G68), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(new_n254), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT12), .B1(new_n271), .B2(G68), .ZN(new_n272));
  OR3_X1    g0072(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(G68), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  OAI211_X1 g0080(.A(G226), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(G232), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT71), .ZN(new_n284));
  OR2_X1    g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT71), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(G232), .A4(G1698), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n282), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G97), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n277), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n267), .B(G274), .C1(G41), .C2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n277), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n294), .B1(new_n297), .B2(G238), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT13), .B1(new_n292), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT13), .ZN(new_n301));
  INV_X1    g0101(.A(new_n291), .ZN(new_n302));
  AOI211_X1 g0102(.A(new_n302), .B(new_n282), .C1(new_n289), .C2(new_n284), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n301), .B(new_n298), .C1(new_n303), .C2(new_n277), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n308), .A3(G169), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n300), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n292), .A2(new_n299), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n275), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n278), .A2(G232), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n287), .B(new_n318), .C1(new_n319), .C2(new_n278), .ZN(new_n320));
  INV_X1    g0120(.A(new_n277), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G107), .C2(new_n287), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n297), .A2(G244), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n293), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n270), .A2(G77), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n231), .A2(G33), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT15), .B(G87), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n271), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(new_n254), .B1(new_n202), .B2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT72), .B1(new_n305), .B2(G200), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT72), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n300), .C2(new_n304), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n313), .A2(new_n315), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n275), .B1(new_n343), .B2(G190), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT74), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n342), .B2(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n317), .B(new_n337), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n278), .A2(G222), .ZN(new_n349));
  INV_X1    g0149(.A(G223), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n287), .B(new_n349), .C1(new_n350), .C2(new_n278), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G77), .B2(new_n287), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT67), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n351), .B(new_n354), .C1(G77), .C2(new_n287), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n321), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n294), .B1(new_n297), .B2(G226), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  INV_X1    g0160(.A(G150), .ZN(new_n361));
  OAI221_X1 g0161(.A(KEYINPUT69), .B1(new_n361), .B2(new_n262), .C1(new_n259), .C2(new_n329), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n329), .B1(new_n257), .B2(new_n258), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n262), .A2(new_n361), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n201), .ZN(new_n367));
  OAI21_X1  g0167(.A(G20), .B1(new_n367), .B2(new_n233), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n362), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n254), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n335), .A2(new_n212), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n270), .A2(G50), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(KEYINPUT9), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT9), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n369), .A2(new_n254), .B1(new_n212), .B2(new_n335), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(new_n372), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT70), .B(new_n360), .C1(new_n374), .C2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n359), .A2(new_n340), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT10), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n373), .A2(KEYINPUT9), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n375), .A3(new_n372), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n379), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n360), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n348), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n285), .A2(new_n231), .A3(new_n286), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n279), .A2(new_n280), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(new_n231), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n261), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n231), .B1(new_n233), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n396), .A4(new_n399), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n254), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n329), .A2(new_n335), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n269), .A2(new_n329), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n350), .A2(new_n278), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n213), .A2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n279), .C2(new_n280), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n321), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n277), .A2(G232), .A3(new_n295), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n415), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT75), .B1(new_n415), .B2(new_n293), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT76), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT76), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n414), .B(new_n420), .C1(new_n416), .C2(new_n417), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G169), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n418), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n311), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n408), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n408), .A2(KEYINPUT18), .A3(new_n424), .A4(new_n426), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n419), .A2(new_n421), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n432), .A2(G200), .B1(G190), .B2(new_n418), .ZN(new_n433));
  XOR2_X1   g0233(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n422), .A2(new_n340), .B1(new_n425), .B2(new_n325), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n408), .A2(new_n437), .B1(KEYINPUT77), .B2(KEYINPUT17), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n429), .A2(new_n430), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n358), .A2(new_n423), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(G179), .B2(new_n358), .ZN(new_n441));
  INV_X1    g0241(.A(new_n373), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n324), .A2(G179), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n336), .A2(new_n328), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n324), .A2(new_n423), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n439), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT78), .B1(new_n389), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n348), .A2(new_n449), .A3(new_n388), .A4(new_n452), .ZN(new_n453));
  OR2_X1    g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n224), .A2(new_n278), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n287), .B(new_n455), .C1(G257), .C2(new_n278), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G294), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n277), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G41), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n267), .B(G45), .C1(new_n459), .C2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  OAI211_X1 g0262(.A(G264), .B(new_n277), .C1(new_n460), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT81), .ZN(new_n466));
  OAI21_X1  g0266(.A(G274), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n467), .A2(new_n468), .A3(new_n460), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n458), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G179), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n423), .B2(new_n470), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n231), .B2(G107), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT23), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT23), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n473), .B(new_n476), .C1(new_n231), .C2(G107), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT85), .B1(new_n478), .B2(G20), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT85), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(new_n231), .A3(G33), .A4(G116), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n475), .A2(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  AOI21_X1  g0283(.A(G20), .B1(new_n285), .B2(new_n286), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G87), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n231), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(KEYINPUT22), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n482), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT24), .B(new_n482), .C1(new_n485), .C2(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(new_n254), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT88), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT25), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n335), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n335), .A2(new_n496), .A3(new_n495), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n494), .A2(KEYINPUT25), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n267), .A2(G33), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n271), .A2(new_n501), .A3(new_n230), .A4(new_n253), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n497), .B(new_n500), .C1(G107), .C2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n492), .A2(new_n493), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n493), .B1(new_n492), .B2(new_n504), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n472), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT89), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT89), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n472), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n492), .A2(new_n504), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n470), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n513), .B(new_n515), .C1(new_n325), .C2(new_n514), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  OAI211_X1 g0317(.A(G257), .B(new_n277), .C1(new_n460), .C2(new_n462), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n224), .B1(new_n285), .B2(new_n286), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g0321(.A(G1698), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(G244), .B1(new_n279), .B2(new_n280), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n521), .B1(G33), .B2(G283), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n278), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n469), .B(new_n519), .C1(new_n526), .C2(new_n321), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n517), .B1(new_n527), .B2(new_n340), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n502), .A2(G97), .ZN(new_n529));
  INV_X1    g0329(.A(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n271), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n392), .B2(new_n394), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT79), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n530), .A2(new_n496), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n390), .A2(new_n391), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n231), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT79), .A3(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n537), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n534), .B1(new_n548), .B2(new_n254), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n527), .A2(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n523), .A2(new_n521), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G283), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n525), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n287), .A2(G250), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n278), .B1(new_n554), .B2(KEYINPUT4), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n321), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n460), .B1(new_n466), .B2(new_n465), .ZN(new_n557));
  INV_X1    g0357(.A(new_n467), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n559), .A3(new_n518), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT82), .A3(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n528), .A2(new_n549), .A3(new_n550), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n423), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n527), .A2(new_n311), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT79), .B1(new_n546), .B2(G107), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n536), .B(new_n496), .C1(new_n544), .C2(new_n545), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n266), .B1(new_n567), .B2(new_n543), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n563), .B(new_n564), .C1(new_n568), .C2(new_n534), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n335), .A2(new_n214), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n266), .A2(G116), .A3(new_n271), .A4(new_n501), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n253), .A2(new_n230), .B1(G20), .B2(new_n214), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n552), .B(new_n231), .C1(G33), .C2(new_n530), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n573), .A2(KEYINPUT20), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT20), .B1(new_n573), .B2(new_n574), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n571), .B(new_n572), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n278), .A2(G257), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G264), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n279), .C2(new_n280), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n321), .C1(G303), .C2(new_n287), .ZN(new_n581));
  OAI211_X1 g0381(.A(G270), .B(new_n277), .C1(new_n460), .C2(new_n462), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n559), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n583), .A3(G169), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n583), .A2(new_n311), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n577), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n577), .A2(new_n583), .A3(KEYINPUT21), .A4(G169), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n231), .B(G68), .C1(new_n279), .C2(new_n280), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n223), .A2(new_n530), .A3(new_n496), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n291), .A2(new_n231), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n332), .A2(KEYINPUT19), .A3(new_n530), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT83), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(KEYINPUT83), .B(new_n591), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n254), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n333), .A2(new_n335), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n319), .A2(new_n278), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n287), .B(new_n604), .C1(G244), .C2(new_n278), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n277), .B1(new_n605), .B2(new_n478), .ZN(new_n606));
  AOI21_X1  g0406(.A(G250), .B1(new_n267), .B2(G45), .ZN(new_n607));
  INV_X1    g0407(.A(G45), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n608), .A2(G1), .A3(G274), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n321), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G190), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n606), .B2(new_n610), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n503), .A2(G87), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n603), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n606), .A2(new_n610), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n423), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n333), .B(KEYINPUT84), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n503), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n601), .A2(new_n602), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n311), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n583), .A2(G200), .ZN(new_n623));
  INV_X1    g0423(.A(new_n577), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n624), .C1(new_n325), .C2(new_n583), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n590), .A2(new_n615), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n570), .A2(new_n626), .ZN(new_n627));
  AND4_X1   g0427(.A1(new_n454), .A2(new_n511), .A3(new_n516), .A4(new_n627), .ZN(G372));
  AND3_X1   g0428(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n613), .A2(new_n601), .A3(new_n614), .A4(new_n602), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n630), .A2(new_n631), .B1(G190), .B2(new_n611), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(new_n516), .A3(new_n569), .A4(new_n562), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n472), .A2(KEYINPUT91), .A3(new_n512), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT91), .B1(new_n472), .B2(new_n512), .ZN(new_n637));
  INV_X1    g0437(.A(new_n590), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n615), .A2(new_n622), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT26), .B1(new_n641), .B2(new_n569), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n633), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n527), .A2(G169), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n560), .A2(G179), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n549), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n646), .A3(new_n622), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n622), .B(new_n642), .C1(new_n647), .C2(KEYINPUT26), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n454), .B1(new_n640), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n429), .A2(new_n430), .ZN(new_n650));
  INV_X1    g0450(.A(new_n317), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n342), .A2(new_n344), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT74), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n448), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n436), .A2(new_n438), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n650), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n380), .A2(KEYINPUT92), .A3(new_n387), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT92), .B1(new_n380), .B2(new_n387), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n443), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n649), .A2(new_n664), .ZN(G369));
  OR2_X1    g0465(.A1(new_n505), .A2(new_n506), .ZN(new_n666));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n267), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n511), .A2(new_n516), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n666), .A2(new_n472), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n674), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n624), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n638), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n590), .A2(new_n625), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n590), .A2(new_n674), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n511), .A2(new_n516), .A3(new_n675), .A4(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n680), .B1(new_n636), .B2(new_n637), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n208), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n593), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n234), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n680), .B1(new_n640), .B2(new_n648), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n635), .B1(new_n511), .B2(new_n590), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n641), .A2(new_n569), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT26), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n629), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(KEYINPUT29), .B(new_n680), .C1(new_n702), .C2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n511), .A2(new_n627), .A3(new_n516), .A4(new_n680), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n458), .A2(new_n464), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n527), .A2(new_n711), .A3(new_n611), .A4(new_n587), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n583), .A2(new_n311), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n514), .A2(new_n560), .A3(new_n616), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(new_n713), .B2(new_n712), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT93), .B1(new_n714), .B2(new_n716), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT31), .B(new_n674), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n712), .A2(new_n713), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n674), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n710), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n709), .B1(G330), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n698), .B1(new_n727), .B2(G1), .ZN(G364));
  OR2_X1    g0528(.A1(new_n684), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n668), .A2(G45), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n694), .A2(G1), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(new_n685), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n230), .B1(G20), .B2(new_n423), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT96), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n231), .A2(new_n325), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n340), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n223), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n231), .A2(G190), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n393), .B(new_n741), .C1(G107), .C2(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT97), .Z(new_n746));
  NOR2_X1   g0546(.A1(G179), .A2(G200), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n231), .B1(new_n747), .B2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G97), .ZN(new_n750));
  INV_X1    g0550(.A(G68), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n311), .A2(new_n340), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n742), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n311), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(KEYINPUT98), .B1(G58), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n738), .A2(new_n752), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n756), .A2(new_n742), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n760), .A2(new_n212), .B1(new_n761), .B2(new_n202), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT98), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n742), .A2(new_n747), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT32), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n746), .A2(new_n759), .A3(new_n764), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n761), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n753), .ZN(new_n772));
  INV_X1    g0572(.A(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(KEYINPUT33), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n765), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G329), .ZN(new_n778));
  INV_X1    g0578(.A(G283), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n776), .B(new_n778), .C1(new_n779), .C2(new_n743), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n771), .B(new_n780), .C1(G294), .C2(new_n749), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n758), .A2(G322), .ZN(new_n782));
  INV_X1    g0582(.A(new_n740), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G303), .ZN(new_n784));
  INV_X1    g0584(.A(new_n760), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n287), .B1(new_n785), .B2(G326), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n781), .A2(new_n782), .A3(new_n784), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n737), .B1(new_n769), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n731), .B(KEYINPUT94), .Z(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT95), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n736), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n248), .A2(G45), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n692), .A2(new_n287), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n608), .B2(new_n235), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n795), .A2(new_n798), .B1(new_n214), .B2(new_n692), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n287), .A2(G355), .A3(new_n208), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n794), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n788), .A2(new_n789), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n792), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n684), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n732), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n726), .A2(G330), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT101), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n446), .A2(new_n674), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n337), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n448), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n656), .A2(new_n680), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n699), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n807), .A2(new_n808), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(new_n731), .C1(new_n816), .C2(new_n809), .ZN(new_n819));
  INV_X1    g0619(.A(new_n791), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n736), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n789), .B1(new_n202), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT99), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n744), .A2(G87), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n824), .B1(new_n779), .B2(new_n753), .C1(new_n770), .C2(new_n765), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n750), .B1(new_n214), .B2(new_n761), .C1(new_n826), .C2(new_n760), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n825), .A2(new_n827), .A3(new_n287), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n496), .B2(new_n740), .C1(new_n829), .C2(new_n757), .ZN(new_n830));
  INV_X1    g0630(.A(new_n761), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G143), .A2(new_n758), .B1(new_n831), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n832), .B1(new_n833), .B2(new_n760), .C1(new_n361), .C2(new_n753), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT34), .Z(new_n835));
  NOR2_X1   g0635(.A1(new_n743), .A2(new_n751), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G50), .B2(new_n783), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n393), .B1(new_n777), .B2(G132), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n749), .A2(G58), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n830), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT100), .Z(new_n842));
  OAI221_X1 g0642(.A(new_n823), .B1(new_n791), .B2(new_n815), .C1(new_n842), .C2(new_n737), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n819), .A2(new_n843), .ZN(G384));
  OAI211_X1 g0644(.A(KEYINPUT31), .B(new_n674), .C1(new_n717), .C2(new_n722), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n710), .A2(new_n725), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n454), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT105), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n317), .B1(new_n346), .B2(new_n347), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n275), .A2(new_n674), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n317), .B(new_n850), .C1(new_n346), .C2(new_n347), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n854), .A2(new_n815), .A3(new_n846), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n650), .A2(new_n658), .ZN(new_n858));
  INV_X1    g0658(.A(new_n672), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n408), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n439), .B2(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n431), .A2(KEYINPUT103), .A3(new_n433), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT103), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n408), .B2(new_n437), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n865), .A2(new_n427), .A3(new_n867), .A4(new_n860), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n431), .A2(new_n433), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT37), .B1(new_n408), .B2(new_n859), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n870), .A2(new_n871), .A3(new_n427), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n862), .A2(new_n864), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n408), .B2(new_n859), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n408), .A2(new_n878), .A3(new_n859), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n858), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n408), .A2(new_n878), .A3(new_n859), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n427), .B(new_n870), .C1(new_n885), .C2(new_n879), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n884), .B(KEYINPUT38), .C1(new_n887), .C2(new_n872), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n857), .B1(new_n877), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n872), .B1(new_n886), .B2(KEYINPUT37), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n882), .B1(new_n650), .B2(new_n658), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n876), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n814), .B1(new_n852), .B2(new_n853), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n846), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n856), .A2(new_n889), .B1(new_n895), .B2(new_n857), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n848), .B(new_n896), .Z(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n888), .A2(new_n892), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n813), .B1(new_n699), .B2(new_n814), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n854), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n899), .A2(new_n901), .B1(new_n650), .B2(new_n859), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT39), .B1(new_n877), .B2(new_n888), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n888), .A2(new_n892), .A3(KEYINPUT39), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n317), .A2(new_n674), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n709), .B1(new_n451), .B2(new_n453), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n664), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n898), .B(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n267), .B2(new_n668), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n214), .B1(new_n542), .B2(KEYINPUT35), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n232), .C1(KEYINPUT35), .C2(new_n542), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT36), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n235), .A2(G77), .A3(new_n397), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n367), .A2(new_n751), .ZN(new_n918));
  OAI211_X1 g0718(.A(G1), .B(new_n667), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT106), .Z(G367));
  OAI211_X1 g0721(.A(new_n562), .B(new_n569), .C1(new_n549), .C2(new_n680), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT107), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n688), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  INV_X1    g0729(.A(new_n511), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n646), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n674), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n603), .A2(new_n614), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n674), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n634), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n629), .A2(new_n933), .A3(new_n674), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR3_X1    g0737(.A1(new_n932), .A2(KEYINPUT43), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n932), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n686), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n924), .B(new_n925), .C1(new_n569), .C2(new_n680), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n938), .A2(new_n686), .A3(new_n945), .A4(new_n942), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT108), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n693), .B(KEYINPUT41), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n946), .A2(new_n690), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n946), .A2(new_n690), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT110), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n946), .A2(KEYINPUT44), .A3(new_n690), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(KEYINPUT110), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n686), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n954), .A2(new_n958), .A3(new_n944), .A4(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n678), .A2(new_n687), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT111), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n688), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n685), .B(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n685), .A2(KEYINPUT112), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n966), .A2(new_n688), .A3(new_n967), .A4(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n970), .A2(new_n727), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT113), .B1(new_n964), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT113), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n962), .A2(new_n973), .A3(new_n976), .A4(new_n963), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n951), .B1(new_n978), .B2(new_n727), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n730), .A2(G1), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n947), .B(new_n949), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n937), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n789), .B1(new_n982), .B2(new_n792), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n793), .B1(new_n208), .B2(new_n333), .C1(new_n243), .C2(new_n797), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n743), .A2(new_n530), .B1(new_n765), .B2(new_n773), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n393), .B1(new_n748), .B2(new_n496), .C1(new_n826), .C2(new_n757), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G283), .C2(new_n831), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n785), .A2(G311), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n783), .A2(G116), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n772), .A2(G294), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n785), .A2(G143), .B1(new_n749), .B2(G68), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n833), .B2(new_n765), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G159), .B2(new_n772), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n744), .A2(G77), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n201), .C2(new_n761), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n287), .B1(new_n757), .B2(new_n361), .C1(new_n247), .C2(new_n740), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI211_X1 g0800(.A(new_n983), .B(new_n984), .C1(new_n737), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n981), .A2(new_n1001), .ZN(G387));
  AND2_X1   g0802(.A1(new_n970), .A2(new_n972), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(new_n727), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n693), .A3(new_n974), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n679), .A2(new_n792), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n783), .A2(G294), .B1(new_n749), .B2(G283), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G322), .A2(new_n785), .B1(new_n772), .B2(G311), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n826), .B2(new_n761), .C1(new_n773), .C2(new_n757), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT115), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT49), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n287), .B1(new_n777), .B2(G326), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n214), .C2(new_n743), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n618), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1018), .A2(new_n748), .B1(new_n766), .B2(new_n760), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n393), .B1(new_n777), .B2(G150), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n202), .B2(new_n740), .C1(new_n530), .C2(new_n743), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT114), .Z(new_n1022));
  AOI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(G50), .C2(new_n758), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n751), .B2(new_n761), .C1(new_n329), .C2(new_n753), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n737), .B1(new_n1017), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n796), .B1(new_n240), .B2(new_n608), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n287), .A2(new_n208), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n695), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n329), .A2(G50), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(G68), .A2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1030), .A2(new_n608), .A3(new_n1031), .A4(new_n695), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n692), .A2(new_n496), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n794), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1025), .A2(new_n789), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1003), .A2(new_n980), .B1(new_n1006), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1005), .A2(new_n1037), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n964), .A2(new_n974), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n978), .A2(new_n1039), .A3(new_n693), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n962), .A2(new_n980), .A3(new_n963), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n793), .B1(new_n530), .B2(new_n208), .C1(new_n251), .C2(new_n797), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n760), .A2(new_n773), .B1(new_n757), .B2(new_n770), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT52), .Z(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G116), .B2(new_n749), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n496), .A2(new_n743), .B1(new_n761), .B2(new_n829), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n287), .B(new_n1046), .C1(G322), .C2(new_n777), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n779), .B2(new_n740), .C1(new_n826), .C2(new_n753), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n748), .A2(new_n202), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G68), .A2(new_n783), .B1(new_n831), .B2(new_n330), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n201), .B2(new_n753), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G143), .C2(new_n777), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n760), .A2(new_n361), .B1(new_n757), .B2(new_n766), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n287), .A3(new_n824), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n789), .B1(new_n1057), .B2(new_n736), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1042), .B(new_n1058), .C1(new_n945), .C2(new_n803), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1040), .A2(new_n1041), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(G390));
  INV_X1    g0861(.A(G125), .ZN(new_n1062));
  INV_X1    g0862(.A(G132), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n287), .B1(new_n765), .B2(new_n1062), .C1(new_n1063), .C2(new_n757), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n783), .A2(G150), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT53), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1064), .B(new_n1066), .C1(G159), .C2(new_n749), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n785), .A2(G128), .B1(new_n744), .B2(new_n367), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(KEYINPUT54), .B(G143), .Z(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n831), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n833), .B2(new_n753), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n741), .A2(new_n836), .A3(new_n1050), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n287), .B1(new_n772), .B2(G107), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G97), .A2(new_n831), .B1(new_n777), .B2(G294), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n214), .B2(new_n757), .C1(new_n779), .C2(new_n760), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n737), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n789), .B(new_n1078), .C1(new_n329), .C2(new_n821), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n906), .B2(new_n791), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n907), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n901), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n903), .B2(new_n905), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n877), .A2(new_n888), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n680), .B(new_n812), .C1(new_n702), .C2(new_n707), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n813), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n854), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1087), .A3(new_n1081), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n726), .A2(G330), .A3(new_n815), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n854), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1083), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n890), .A2(new_n891), .A3(new_n876), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n876), .B2(new_n875), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n904), .B1(new_n1093), .B2(KEYINPUT39), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n907), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1094), .A2(new_n1082), .B1(new_n1095), .B2(new_n1087), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n894), .A2(G330), .A3(new_n846), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n980), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1080), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n846), .C1(new_n451), .C2(new_n453), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1101), .A2(new_n664), .A3(new_n909), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n850), .B1(new_n655), .B2(new_n317), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n853), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n815), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n846), .A2(G330), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1105), .A2(new_n1106), .B1(new_n1089), .B2(new_n854), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n900), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n854), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n846), .A2(KEYINPUT116), .A3(G330), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n815), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT116), .B1(new_n846), .B2(G330), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1086), .B1(new_n1089), .B2(new_n854), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1102), .A2(new_n1116), .A3(KEYINPUT117), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n900), .A2(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1101), .A2(new_n664), .A3(new_n909), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1097), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1096), .B2(new_n1090), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n694), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1098), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1100), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G378));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1120), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1084), .A2(KEYINPUT40), .A3(new_n846), .A4(new_n894), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n857), .B1(new_n855), .B2(new_n899), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(G330), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n373), .A2(new_n859), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT118), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n663), .B2(new_n444), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n661), .A2(new_n662), .A3(new_n443), .A4(new_n1137), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n662), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n380), .A2(KEYINPUT92), .A3(new_n387), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n444), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n663), .A2(new_n444), .A3(new_n1138), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n1135), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1133), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n1131), .A3(new_n1132), .A4(G330), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1150), .A2(new_n908), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n908), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1129), .B1(new_n1130), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1148), .B1(new_n896), .B2(G330), .ZN(new_n1156));
  AND4_X1   g0956(.A1(G330), .A2(new_n1148), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1094), .A2(new_n1081), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(new_n902), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1150), .A2(new_n908), .A3(new_n1151), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1098), .B1(new_n1121), .B2(new_n1117), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(KEYINPUT57), .C1(new_n1162), .C2(new_n1120), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1155), .A2(new_n693), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1149), .A2(new_n820), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n821), .A2(new_n201), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n459), .B1(new_n748), .B2(new_n751), .C1(new_n202), .C2(new_n740), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G58), .A2(new_n744), .B1(new_n777), .B2(G283), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n393), .C1(new_n530), .C2(new_n753), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1167), .B(new_n1169), .C1(G116), .C2(new_n785), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n496), .B2(new_n757), .C1(new_n1018), .C2(new_n761), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n212), .B1(new_n279), .B2(G41), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G128), .A2(new_n758), .B1(new_n831), .B2(G137), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n783), .A2(new_n1070), .B1(new_n749), .B2(G150), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n1062), .C2(new_n760), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G132), .B2(new_n772), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G41), .B1(new_n777), .B2(G124), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n256), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G159), .B2(new_n744), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1178), .B2(new_n1177), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1172), .A2(new_n1173), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n731), .B1(new_n1184), .B2(new_n736), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1165), .A2(new_n1166), .A3(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT119), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n1099), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1117), .A2(new_n1121), .A3(new_n950), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1109), .A2(new_n820), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n785), .A2(G132), .B1(new_n831), .B2(G150), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n833), .B2(new_n757), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G159), .A2(new_n783), .B1(new_n777), .B2(G128), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT121), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n772), .C2(new_n1070), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1198), .B(new_n287), .C1(new_n212), .C2(new_n748), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G58), .B2(new_n744), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n618), .A2(new_n749), .B1(G97), .B2(new_n783), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n829), .B2(new_n760), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G116), .B2(new_n772), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n996), .B1(new_n496), .B2(new_n761), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n287), .B(new_n1204), .C1(G303), .C2(new_n777), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n779), .C2(new_n757), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT120), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n736), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n789), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n821), .A2(new_n751), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT122), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1116), .A2(new_n980), .B1(new_n1193), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1192), .A2(new_n1213), .ZN(G381));
  NAND3_X1  g1014(.A1(new_n981), .A2(new_n1060), .A3(new_n1001), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G375), .A2(G378), .ZN(new_n1217));
  INV_X1    g1017(.A(G381), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(G407));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n673), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(G213), .A3(new_n1221), .ZN(G409));
  XNOR2_X1  g1022(.A(G393), .B(new_n805), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1060), .B1(new_n981), .B2(new_n1001), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1216), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(G387), .A2(G390), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1223), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1215), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1127), .B1(new_n1164), .B2(new_n1189), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1186), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT123), .B1(new_n1188), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n980), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1186), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1161), .B(new_n950), .C1(new_n1162), .C2(new_n1120), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1232), .A2(new_n1127), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n673), .A2(G213), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1230), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1117), .A2(new_n1121), .A3(KEYINPUT60), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(KEYINPUT124), .A3(new_n1191), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT124), .B1(new_n1242), .B2(new_n1191), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n693), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1213), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1191), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1246), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1242), .A2(KEYINPUT124), .A3(new_n1191), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(G384), .A3(new_n1213), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1249), .A2(KEYINPUT125), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1255), .A2(G384), .A3(new_n1213), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G384), .B1(new_n1255), .B2(new_n1213), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1240), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1240), .A2(new_n1261), .A3(new_n1264), .A4(new_n1257), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n673), .A2(G213), .A3(G2897), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1261), .A2(new_n1268), .A3(new_n1257), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1270), .A2(new_n1268), .B1(new_n1230), .B2(new_n1239), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1229), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1268), .B1(new_n1249), .B2(new_n1256), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1240), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1261), .A2(new_n1268), .A3(new_n1257), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1240), .A2(new_n1261), .A3(KEYINPUT63), .A4(new_n1257), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1262), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1274), .A2(new_n1278), .A3(new_n1279), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1273), .A2(new_n1282), .ZN(G405));
  INV_X1    g1083(.A(KEYINPUT127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1229), .A2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1217), .A2(new_n1230), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1217), .A2(new_n1230), .B1(new_n1260), .B2(new_n1259), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1225), .A2(new_n1228), .A3(KEYINPUT127), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1285), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n1288), .A4(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(G402));
endmodule


