

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793;

  XNOR2_X1 U374 ( .A(n604), .B(KEYINPUT1), .ZN(n644) );
  NAND2_X1 U375 ( .A1(n706), .A2(n370), .ZN(n369) );
  NAND2_X1 U376 ( .A1(n619), .A2(n710), .ZN(n596) );
  NOR2_X2 U377 ( .A1(n470), .A2(n579), .ZN(n531) );
  AND2_X2 U378 ( .A1(n419), .A2(n417), .ZN(n416) );
  NOR2_X2 U379 ( .A1(n791), .A2(n793), .ZN(n454) );
  XNOR2_X2 U380 ( .A(n639), .B(n638), .ZN(n791) );
  NAND2_X2 U381 ( .A1(n416), .A2(n412), .ZN(n674) );
  NAND2_X2 U382 ( .A1(n563), .A2(n355), .ZN(n564) );
  OR2_X2 U383 ( .A1(n664), .A2(G902), .ZN(n502) );
  AND2_X2 U384 ( .A1(n592), .A2(n603), .ZN(n593) );
  INV_X1 U385 ( .A(KEYINPUT92), .ZN(n385) );
  INV_X1 U386 ( .A(KEYINPUT64), .ZN(n372) );
  XNOR2_X1 U387 ( .A(n386), .B(n385), .ZN(n384) );
  NOR2_X1 U388 ( .A1(n440), .A2(n576), .ZN(n684) );
  NOR2_X1 U389 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U390 ( .A1(n606), .A2(n528), .ZN(n530) );
  NAND2_X2 U391 ( .A1(n707), .A2(n628), .ZN(n581) );
  XNOR2_X1 U392 ( .A(n484), .B(n483), .ZN(n723) );
  AND2_X1 U393 ( .A1(n383), .A2(n382), .ZN(n381) );
  XOR2_X1 U394 ( .A(n664), .B(KEYINPUT62), .Z(n478) );
  XNOR2_X1 U395 ( .A(n397), .B(n511), .ZN(n664) );
  XNOR2_X1 U396 ( .A(n505), .B(n493), .ZN(n497) );
  XNOR2_X1 U397 ( .A(n372), .B(G953), .ZN(n506) );
  INV_X1 U398 ( .A(KEYINPUT119), .ZN(n438) );
  BUF_X1 U399 ( .A(G128), .Z(n407) );
  BUF_X1 U400 ( .A(n470), .Z(n351) );
  XNOR2_X1 U401 ( .A(n455), .B(n360), .ZN(n470) );
  NOR2_X1 U402 ( .A1(G953), .A2(n752), .ZN(n753) );
  XNOR2_X1 U403 ( .A(n439), .B(n438), .ZN(n752) );
  NAND2_X1 U404 ( .A1(n389), .A2(n384), .ZN(n352) );
  NAND2_X1 U405 ( .A1(n389), .A2(n384), .ZN(n428) );
  AND2_X1 U406 ( .A1(n392), .A2(n390), .ZN(n389) );
  AND2_X1 U407 ( .A1(n769), .A2(n584), .ZN(n655) );
  NAND2_X1 U408 ( .A1(n430), .A2(KEYINPUT36), .ZN(n420) );
  NAND2_X2 U409 ( .A1(n381), .A2(n377), .ZN(n604) );
  NAND2_X1 U410 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U411 ( .A(G472), .ZN(n461) );
  XNOR2_X1 U412 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U413 ( .A(KEYINPUT25), .ZN(n481) );
  AND2_X1 U414 ( .A1(n466), .A2(n465), .ZN(n464) );
  INV_X1 U415 ( .A(KEYINPUT74), .ZN(n462) );
  NAND2_X1 U416 ( .A1(n437), .A2(n436), .ZN(n572) );
  XNOR2_X1 U417 ( .A(n391), .B(n429), .ZN(n390) );
  INV_X1 U418 ( .A(KEYINPUT65), .ZN(n429) );
  NAND2_X1 U419 ( .A1(n572), .A2(KEYINPUT44), .ZN(n391) );
  XNOR2_X1 U420 ( .A(n513), .B(G122), .ZN(n534) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n513) );
  INV_X1 U422 ( .A(G478), .ZN(n371) );
  XNOR2_X1 U423 ( .A(G131), .B(G134), .ZN(n493) );
  NOR2_X2 U424 ( .A1(G953), .A2(G237), .ZN(n539) );
  XNOR2_X1 U425 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U426 ( .A(G146), .B(G137), .ZN(n375) );
  XNOR2_X1 U427 ( .A(n373), .B(G116), .ZN(n376) );
  INV_X1 U428 ( .A(KEYINPUT5), .ZN(n373) );
  XNOR2_X1 U429 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n498) );
  XNOR2_X1 U430 ( .A(n452), .B(n451), .ZN(n532) );
  INV_X1 U431 ( .A(KEYINPUT8), .ZN(n451) );
  NAND2_X1 U432 ( .A1(n506), .A2(G234), .ZN(n452) );
  XNOR2_X1 U433 ( .A(n534), .B(n533), .ZN(n366) );
  XOR2_X1 U434 ( .A(G134), .B(KEYINPUT105), .Z(n533) );
  NAND2_X1 U435 ( .A1(n532), .A2(G217), .ZN(n367) );
  AND2_X1 U436 ( .A1(n432), .A2(n445), .ZN(n431) );
  NAND2_X1 U437 ( .A1(n433), .A2(KEYINPUT36), .ZN(n432) );
  INV_X1 U438 ( .A(KEYINPUT111), .ZN(n414) );
  NAND2_X1 U439 ( .A1(n357), .A2(n566), .ZN(n475) );
  NOR2_X1 U440 ( .A1(n402), .A2(n761), .ZN(n401) );
  NAND2_X1 U441 ( .A1(n410), .A2(n361), .ZN(n400) );
  NOR2_X1 U442 ( .A1(n447), .A2(G210), .ZN(n402) );
  XOR2_X1 U443 ( .A(n642), .B(KEYINPUT48), .Z(n476) );
  NAND2_X1 U444 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U445 ( .A1(n684), .A2(n356), .ZN(n388) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n522) );
  OR2_X1 U447 ( .A1(G237), .A2(G902), .ZN(n520) );
  INV_X1 U448 ( .A(G469), .ZN(n380) );
  NAND2_X1 U449 ( .A1(G902), .A2(G469), .ZN(n382) );
  XNOR2_X1 U450 ( .A(G902), .B(KEYINPUT15), .ZN(n658) );
  XNOR2_X1 U451 ( .A(G113), .B(KEYINPUT103), .ZN(n547) );
  XNOR2_X1 U452 ( .A(G131), .B(KEYINPUT12), .ZN(n548) );
  XNOR2_X1 U453 ( .A(G140), .B(KEYINPUT101), .ZN(n541) );
  XNOR2_X1 U454 ( .A(n540), .B(KEYINPUT102), .ZN(n542) );
  XNOR2_X1 U455 ( .A(G104), .B(KEYINPUT11), .ZN(n545) );
  XNOR2_X1 U456 ( .A(G107), .B(G146), .ZN(n489) );
  XNOR2_X1 U457 ( .A(G104), .B(KEYINPUT97), .ZN(n492) );
  XNOR2_X1 U458 ( .A(G137), .B(G140), .ZN(n408) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT95), .Z(n508) );
  INV_X1 U460 ( .A(n597), .ZN(n433) );
  INV_X1 U461 ( .A(KEYINPUT80), .ZN(n457) );
  NOR2_X1 U462 ( .A1(n614), .A2(n615), .ZN(n616) );
  XNOR2_X1 U463 ( .A(n530), .B(n529), .ZN(n561) );
  XNOR2_X1 U464 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n529) );
  OR2_X1 U465 ( .A1(n675), .A2(G902), .ZN(n556) );
  XNOR2_X1 U466 ( .A(G137), .B(G140), .ZN(n494) );
  XNOR2_X1 U467 ( .A(n425), .B(G128), .ZN(n424) );
  INV_X1 U468 ( .A(G119), .ZN(n425) );
  XNOR2_X1 U469 ( .A(n473), .B(KEYINPUT24), .ZN(n472) );
  XNOR2_X1 U470 ( .A(KEYINPUT23), .B(G110), .ZN(n473) );
  XNOR2_X1 U471 ( .A(n427), .B(n426), .ZN(n605) );
  XNOR2_X1 U472 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n426) );
  NAND2_X1 U473 ( .A1(n460), .A2(n603), .ZN(n427) );
  INV_X1 U474 ( .A(n456), .ZN(n460) );
  BUF_X1 U475 ( .A(n727), .Z(n456) );
  XNOR2_X1 U476 ( .A(n497), .B(n396), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n374), .B(n496), .ZN(n396) );
  BUF_X1 U478 ( .A(n506), .Z(n786) );
  XNOR2_X1 U479 ( .A(n367), .B(n366), .ZN(n368) );
  NAND2_X1 U480 ( .A1(n750), .A2(n751), .ZN(n439) );
  NAND2_X1 U481 ( .A1(n415), .A2(n413), .ZN(n412) );
  INV_X1 U482 ( .A(n421), .ZN(n415) );
  INV_X1 U483 ( .A(KEYINPUT66), .ZN(n567) );
  NOR2_X1 U484 ( .A1(n369), .A2(n460), .ZN(n685) );
  INV_X1 U485 ( .A(KEYINPUT120), .ZN(n442) );
  INV_X1 U486 ( .A(KEYINPUT56), .ZN(n444) );
  NAND2_X1 U487 ( .A1(n398), .A2(n354), .ZN(n395) );
  NOR2_X1 U488 ( .A1(n456), .A2(n459), .ZN(n353) );
  AND2_X1 U489 ( .A1(n400), .A2(n401), .ZN(n354) );
  AND2_X1 U490 ( .A1(n590), .A2(n562), .ZN(n355) );
  AND2_X1 U491 ( .A1(n583), .A2(n582), .ZN(n356) );
  XNOR2_X1 U492 ( .A(KEYINPUT107), .B(n565), .ZN(n357) );
  AND2_X1 U493 ( .A1(n704), .A2(n652), .ZN(n358) );
  NOR2_X1 U494 ( .A1(n351), .A2(n740), .ZN(n359) );
  INV_X1 U495 ( .A(G902), .ZN(n379) );
  INV_X1 U496 ( .A(n710), .ZN(n459) );
  XOR2_X1 U497 ( .A(KEYINPUT94), .B(KEYINPUT33), .Z(n360) );
  AND2_X1 U498 ( .A1(n447), .A2(G210), .ZN(n361) );
  XNOR2_X1 U499 ( .A(n567), .B(KEYINPUT32), .ZN(n474) );
  XOR2_X1 U500 ( .A(n679), .B(n678), .Z(n362) );
  XNOR2_X1 U501 ( .A(KEYINPUT59), .B(n675), .ZN(n363) );
  XNOR2_X1 U502 ( .A(n666), .B(KEYINPUT96), .ZN(n761) );
  INV_X1 U503 ( .A(n761), .ZN(n446) );
  XOR2_X1 U504 ( .A(n659), .B(KEYINPUT67), .Z(n364) );
  XNOR2_X1 U505 ( .A(n677), .B(KEYINPUT68), .ZN(n365) );
  XNOR2_X1 U506 ( .A(n368), .B(n537), .ZN(n754) );
  NOR2_X1 U507 ( .A1(n706), .A2(n707), .ZN(n621) );
  INV_X1 U508 ( .A(n369), .ZN(n651) );
  NOR2_X1 U509 ( .A1(n629), .A2(n370), .ZN(n630) );
  INV_X1 U510 ( .A(n707), .ZN(n370) );
  XNOR2_X2 U511 ( .A(n538), .B(n371), .ZN(n707) );
  OR2_X1 U512 ( .A1(n679), .A2(n378), .ZN(n377) );
  NAND2_X1 U513 ( .A1(n679), .A2(G469), .ZN(n383) );
  XNOR2_X1 U514 ( .A(n495), .B(n780), .ZN(n679) );
  NAND2_X1 U515 ( .A1(n406), .A2(KEYINPUT44), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n394), .A2(n393), .ZN(n392) );
  XNOR2_X1 U517 ( .A(n572), .B(KEYINPUT93), .ZN(n393) );
  XNOR2_X1 U518 ( .A(n560), .B(n422), .ZN(n394) );
  XNOR2_X1 U519 ( .A(n395), .B(n444), .ZN(G51) );
  XNOR2_X2 U520 ( .A(n535), .B(n469), .ZN(n505) );
  NAND2_X1 U521 ( .A1(n399), .A2(n683), .ZN(n398) );
  INV_X1 U522 ( .A(n410), .ZN(n399) );
  XNOR2_X1 U523 ( .A(n352), .B(KEYINPUT45), .ZN(n403) );
  XNOR2_X1 U524 ( .A(n428), .B(KEYINPUT45), .ZN(n769) );
  XNOR2_X1 U525 ( .A(n564), .B(KEYINPUT22), .ZN(n404) );
  XNOR2_X1 U526 ( .A(n564), .B(KEYINPUT22), .ZN(n568) );
  BUF_X1 U527 ( .A(n754), .Z(n405) );
  XNOR2_X1 U528 ( .A(n559), .B(KEYINPUT35), .ZN(n406) );
  XNOR2_X1 U529 ( .A(n559), .B(KEYINPUT35), .ZN(n790) );
  XNOR2_X1 U530 ( .A(n497), .B(n408), .ZN(n780) );
  XNOR2_X1 U531 ( .A(n503), .B(KEYINPUT10), .ZN(n778) );
  XNOR2_X1 U532 ( .A(n437), .B(G119), .ZN(G21) );
  XNOR2_X1 U533 ( .A(n449), .B(n491), .ZN(n495) );
  XNOR2_X1 U534 ( .A(n490), .B(n514), .ZN(n449) );
  BUF_X1 U535 ( .A(n723), .Z(n440) );
  XOR2_X1 U536 ( .A(G143), .B(n407), .Z(n409) );
  AND2_X1 U537 ( .A1(n784), .A2(n657), .ZN(n747) );
  AND2_X2 U538 ( .A1(n663), .A2(n743), .ZN(n410) );
  AND2_X2 U539 ( .A1(n663), .A2(n743), .ZN(n757) );
  BUF_X1 U540 ( .A(n661), .Z(n784) );
  XNOR2_X2 U541 ( .A(n581), .B(n580), .ZN(n411) );
  XNOR2_X1 U542 ( .A(n581), .B(n580), .ZN(n697) );
  NOR2_X1 U543 ( .A1(n404), .A2(n570), .ZN(n571) );
  AND2_X1 U544 ( .A1(n420), .A2(n414), .ZN(n413) );
  NAND2_X1 U545 ( .A1(n418), .A2(KEYINPUT111), .ZN(n417) );
  INV_X1 U546 ( .A(n420), .ZN(n418) );
  NAND2_X1 U547 ( .A1(n421), .A2(KEYINPUT111), .ZN(n419) );
  XNOR2_X1 U548 ( .A(n674), .B(n468), .ZN(n467) );
  NAND2_X1 U549 ( .A1(n434), .A2(n431), .ZN(n421) );
  INV_X1 U550 ( .A(KEYINPUT71), .ZN(n422) );
  XNOR2_X1 U551 ( .A(n423), .B(n472), .ZN(n471) );
  XNOR2_X1 U552 ( .A(n424), .B(n494), .ZN(n423) );
  XNOR2_X2 U553 ( .A(n453), .B(n474), .ZN(n437) );
  INV_X1 U554 ( .A(n598), .ZN(n430) );
  NAND2_X1 U555 ( .A1(n598), .A2(n435), .ZN(n434) );
  AND2_X1 U556 ( .A1(n597), .A2(n599), .ZN(n435) );
  INV_X1 U557 ( .A(n571), .ZN(n436) );
  NAND2_X1 U558 ( .A1(n757), .A2(G475), .ZN(n676) );
  XNOR2_X1 U559 ( .A(n441), .B(n365), .ZN(G60) );
  NAND2_X1 U560 ( .A1(n450), .A2(n446), .ZN(n441) );
  NAND2_X1 U561 ( .A1(n653), .A2(n358), .ZN(n661) );
  XNOR2_X1 U562 ( .A(n443), .B(n442), .ZN(G54) );
  NAND2_X1 U563 ( .A1(n448), .A2(n446), .ZN(n443) );
  BUF_X1 U564 ( .A(n644), .Z(n445) );
  INV_X1 U565 ( .A(n683), .ZN(n447) );
  XNOR2_X1 U566 ( .A(n680), .B(n362), .ZN(n448) );
  NAND2_X1 U567 ( .A1(n660), .A2(n364), .ZN(n663) );
  XNOR2_X1 U568 ( .A(n676), .B(n363), .ZN(n450) );
  NAND2_X1 U569 ( .A1(n577), .A2(n460), .ZN(n731) );
  NAND2_X1 U570 ( .A1(n593), .A2(n411), .ZN(n595) );
  NOR2_X2 U571 ( .A1(n404), .A2(n475), .ZN(n453) );
  XNOR2_X1 U572 ( .A(n471), .B(n778), .ZN(n479) );
  XNOR2_X1 U573 ( .A(n454), .B(KEYINPUT46), .ZN(n640) );
  XNOR2_X1 U574 ( .A(n643), .B(n476), .ZN(n653) );
  NAND2_X1 U575 ( .A1(n650), .A2(n411), .ZN(n639) );
  XNOR2_X2 U576 ( .A(n637), .B(KEYINPUT39), .ZN(n650) );
  BUF_X2 U577 ( .A(n561), .Z(n579) );
  INV_X1 U578 ( .A(n701), .ZN(n698) );
  XNOR2_X1 U579 ( .A(n578), .B(KEYINPUT31), .ZN(n701) );
  NAND2_X1 U580 ( .A1(n577), .A2(n592), .ZN(n455) );
  INV_X1 U581 ( .A(n628), .ZN(n706) );
  XNOR2_X2 U582 ( .A(n556), .B(n555), .ZN(n628) );
  XNOR2_X2 U583 ( .A(n458), .B(n457), .ZN(n577) );
  NAND2_X1 U584 ( .A1(n718), .A2(n644), .ZN(n458) );
  XNOR2_X2 U585 ( .A(n502), .B(n461), .ZN(n727) );
  XNOR2_X1 U586 ( .A(n463), .B(n462), .ZN(n641) );
  NAND2_X1 U587 ( .A1(n467), .A2(n464), .ZN(n463) );
  NAND2_X1 U588 ( .A1(n611), .A2(n610), .ZN(n465) );
  NOR2_X1 U589 ( .A1(n626), .A2(n625), .ZN(n466) );
  INV_X1 U590 ( .A(KEYINPUT90), .ZN(n468) );
  XNOR2_X2 U591 ( .A(KEYINPUT73), .B(KEYINPUT4), .ZN(n469) );
  XNOR2_X2 U592 ( .A(G143), .B(G128), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n717), .A2(n351), .ZN(n736) );
  XNOR2_X2 U594 ( .A(G146), .B(G125), .ZN(n503) );
  AND2_X1 U595 ( .A1(n532), .A2(G221), .ZN(n477) );
  XNOR2_X1 U596 ( .A(n500), .B(n489), .ZN(n490) );
  INV_X1 U597 ( .A(n596), .ZN(n597) );
  XNOR2_X1 U598 ( .A(n479), .B(n477), .ZN(n758) );
  NOR2_X1 U599 ( .A1(n758), .A2(G902), .ZN(n484) );
  NAND2_X1 U600 ( .A1(n658), .A2(G234), .ZN(n480) );
  XNOR2_X1 U601 ( .A(n480), .B(KEYINPUT20), .ZN(n485) );
  NAND2_X1 U602 ( .A1(G217), .A2(n485), .ZN(n482) );
  NAND2_X1 U603 ( .A1(G221), .A2(n485), .ZN(n486) );
  XNOR2_X1 U604 ( .A(KEYINPUT21), .B(n486), .ZN(n724) );
  NOR2_X2 U605 ( .A1(n723), .A2(n724), .ZN(n487) );
  XNOR2_X2 U606 ( .A(n487), .B(KEYINPUT72), .ZN(n718) );
  NAND2_X1 U607 ( .A1(G227), .A2(n786), .ZN(n491) );
  INV_X1 U608 ( .A(KEYINPUT70), .ZN(n488) );
  XNOR2_X1 U609 ( .A(n488), .B(G101), .ZN(n500) );
  XNOR2_X1 U610 ( .A(n492), .B(G110), .ZN(n514) );
  NAND2_X1 U611 ( .A1(n539), .A2(G210), .ZN(n496) );
  XOR2_X1 U612 ( .A(G113), .B(G119), .Z(n499) );
  XNOR2_X1 U613 ( .A(n499), .B(n498), .ZN(n764) );
  INV_X1 U614 ( .A(n500), .ZN(n501) );
  XNOR2_X1 U615 ( .A(n764), .B(n501), .ZN(n511) );
  XNOR2_X2 U616 ( .A(n727), .B(KEYINPUT6), .ZN(n592) );
  XNOR2_X1 U617 ( .A(n503), .B(KEYINPUT18), .ZN(n504) );
  XNOR2_X1 U618 ( .A(n504), .B(n505), .ZN(n510) );
  NAND2_X1 U619 ( .A1(G224), .A2(n506), .ZN(n507) );
  XNOR2_X1 U620 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n512), .B(n511), .ZN(n517) );
  XOR2_X1 U623 ( .A(n534), .B(KEYINPUT16), .Z(n516) );
  XNOR2_X1 U624 ( .A(n514), .B(KEYINPUT76), .ZN(n515) );
  XNOR2_X1 U625 ( .A(n516), .B(n515), .ZN(n763) );
  XNOR2_X1 U626 ( .A(n517), .B(n763), .ZN(n681) );
  NAND2_X1 U627 ( .A1(n681), .A2(n658), .ZN(n519) );
  AND2_X1 U628 ( .A1(G210), .A2(n520), .ZN(n518) );
  XNOR2_X2 U629 ( .A(n519), .B(n518), .ZN(n619) );
  NAND2_X1 U630 ( .A1(G214), .A2(n520), .ZN(n710) );
  INV_X1 U631 ( .A(KEYINPUT19), .ZN(n521) );
  XNOR2_X2 U632 ( .A(n596), .B(n521), .ZN(n606) );
  XNOR2_X1 U633 ( .A(n522), .B(KEYINPUT98), .ZN(n523) );
  XNOR2_X1 U634 ( .A(KEYINPUT14), .B(n523), .ZN(n525) );
  NAND2_X1 U635 ( .A1(n525), .A2(G952), .ZN(n524) );
  XOR2_X1 U636 ( .A(KEYINPUT99), .B(n524), .Z(n739) );
  NOR2_X1 U637 ( .A1(G953), .A2(n739), .ZN(n589) );
  AND2_X1 U638 ( .A1(n525), .A2(G902), .ZN(n586) );
  INV_X1 U639 ( .A(G953), .ZN(n770) );
  NOR2_X1 U640 ( .A1(G898), .A2(n770), .ZN(n767) );
  NAND2_X1 U641 ( .A1(n586), .A2(n767), .ZN(n526) );
  XOR2_X1 U642 ( .A(KEYINPUT100), .B(n526), .Z(n527) );
  NOR2_X1 U643 ( .A1(n589), .A2(n527), .ZN(n528) );
  XNOR2_X1 U644 ( .A(n531), .B(KEYINPUT34), .ZN(n558) );
  XNOR2_X1 U645 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n409), .B(n536), .ZN(n537) );
  NAND2_X1 U647 ( .A1(n754), .A2(n379), .ZN(n538) );
  NAND2_X1 U648 ( .A1(n539), .A2(G214), .ZN(n540) );
  XNOR2_X1 U649 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U650 ( .A(n543), .B(n778), .ZN(n552) );
  INV_X1 U651 ( .A(G143), .ZN(n544) );
  XNOR2_X1 U652 ( .A(n544), .B(G122), .ZN(n546) );
  XNOR2_X1 U653 ( .A(n546), .B(n545), .ZN(n550) );
  XNOR2_X1 U654 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U655 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U656 ( .A(n552), .B(n551), .ZN(n675) );
  XNOR2_X1 U657 ( .A(KEYINPUT13), .B(G475), .ZN(n554) );
  INV_X1 U658 ( .A(KEYINPUT104), .ZN(n553) );
  XNOR2_X1 U659 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U660 ( .A(KEYINPUT83), .B(n621), .Z(n557) );
  NAND2_X1 U661 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X2 U662 ( .A1(n790), .A2(KEYINPUT44), .ZN(n560) );
  INV_X1 U663 ( .A(n561), .ZN(n563) );
  INV_X1 U664 ( .A(n724), .ZN(n590) );
  AND2_X1 U665 ( .A1(n707), .A2(n706), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n440), .A2(n644), .ZN(n565) );
  XOR2_X1 U667 ( .A(KEYINPUT84), .B(n592), .Z(n566) );
  NAND2_X1 U668 ( .A1(n440), .A2(n456), .ZN(n569) );
  OR2_X1 U669 ( .A1(n569), .A2(n445), .ZN(n570) );
  INV_X1 U670 ( .A(n445), .ZN(n719) );
  INV_X1 U671 ( .A(n592), .ZN(n573) );
  NAND2_X1 U672 ( .A1(n719), .A2(n573), .ZN(n574) );
  NOR2_X1 U673 ( .A1(n568), .A2(n574), .ZN(n575) );
  XNOR2_X1 U674 ( .A(n575), .B(KEYINPUT91), .ZN(n576) );
  NOR2_X1 U675 ( .A1(n579), .A2(n731), .ZN(n578) );
  NAND2_X1 U676 ( .A1(n718), .A2(n604), .ZN(n614) );
  NOR2_X1 U677 ( .A1(n579), .A2(n614), .ZN(n686) );
  NAND2_X1 U678 ( .A1(n686), .A2(n456), .ZN(n670) );
  NAND2_X1 U679 ( .A1(n701), .A2(n670), .ZN(n583) );
  INV_X1 U680 ( .A(KEYINPUT106), .ZN(n580) );
  INV_X1 U681 ( .A(n697), .ZN(n669) );
  NAND2_X1 U682 ( .A1(n669), .A2(n369), .ZN(n712) );
  XNOR2_X1 U683 ( .A(n712), .B(KEYINPUT85), .ZN(n600) );
  INV_X1 U684 ( .A(n600), .ZN(n582) );
  INV_X1 U685 ( .A(n658), .ZN(n584) );
  INV_X1 U686 ( .A(n786), .ZN(n585) );
  NAND2_X1 U687 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U688 ( .A1(G900), .A2(n587), .ZN(n588) );
  OR2_X1 U689 ( .A1(n589), .A2(n588), .ZN(n613) );
  AND2_X1 U690 ( .A1(n613), .A2(n590), .ZN(n591) );
  AND2_X1 U691 ( .A1(n723), .A2(n591), .ZN(n603) );
  INV_X1 U692 ( .A(KEYINPUT108), .ZN(n594) );
  XNOR2_X2 U693 ( .A(n595), .B(n594), .ZN(n646) );
  XNOR2_X1 U694 ( .A(n646), .B(KEYINPUT110), .ZN(n598) );
  INV_X1 U695 ( .A(KEYINPUT36), .ZN(n599) );
  NOR2_X1 U696 ( .A1(KEYINPUT47), .A2(n600), .ZN(n601) );
  XOR2_X1 U697 ( .A(KEYINPUT78), .B(n601), .Z(n612) );
  INV_X1 U698 ( .A(n612), .ZN(n602) );
  INV_X1 U699 ( .A(KEYINPUT77), .ZN(n608) );
  NAND2_X1 U700 ( .A1(n602), .A2(n608), .ZN(n607) );
  NAND2_X1 U701 ( .A1(n605), .A2(n604), .ZN(n632) );
  NOR2_X1 U702 ( .A1(n632), .A2(n606), .ZN(n690) );
  NAND2_X1 U703 ( .A1(n607), .A2(n690), .ZN(n611) );
  INV_X1 U704 ( .A(KEYINPUT47), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n623), .A2(n608), .ZN(n609) );
  OR2_X1 U706 ( .A1(n690), .A2(n609), .ZN(n610) );
  AND2_X1 U707 ( .A1(n612), .A2(KEYINPUT77), .ZN(n626) );
  INV_X1 U708 ( .A(n613), .ZN(n615) );
  XNOR2_X1 U709 ( .A(KEYINPUT82), .B(n616), .ZN(n618) );
  XNOR2_X1 U710 ( .A(n353), .B(KEYINPUT30), .ZN(n617) );
  NAND2_X1 U711 ( .A1(n618), .A2(n617), .ZN(n635) );
  BUF_X1 U712 ( .A(n619), .Z(n620) );
  NAND2_X1 U713 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U714 ( .A1(n635), .A2(n622), .ZN(n696) );
  NOR2_X1 U715 ( .A1(n712), .A2(n623), .ZN(n624) );
  OR2_X1 U716 ( .A1(n696), .A2(n624), .ZN(n625) );
  XOR2_X1 U717 ( .A(KEYINPUT79), .B(KEYINPUT38), .Z(n627) );
  XOR2_X1 U718 ( .A(n620), .B(n627), .Z(n711) );
  OR2_X1 U719 ( .A1(n628), .A2(n459), .ZN(n629) );
  AND2_X1 U720 ( .A1(n711), .A2(n630), .ZN(n631) );
  XNOR2_X1 U721 ( .A(n631), .B(KEYINPUT41), .ZN(n740) );
  NOR2_X1 U722 ( .A1(n740), .A2(n632), .ZN(n633) );
  XNOR2_X1 U723 ( .A(n633), .B(KEYINPUT42), .ZN(n793) );
  INV_X1 U724 ( .A(n711), .ZN(n634) );
  INV_X1 U725 ( .A(n636), .ZN(n637) );
  INV_X1 U726 ( .A(KEYINPUT40), .ZN(n638) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n643) );
  INV_X1 U728 ( .A(KEYINPUT89), .ZN(n642) );
  NOR2_X1 U729 ( .A1(n445), .A2(n459), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n647), .B(KEYINPUT43), .ZN(n649) );
  INV_X1 U732 ( .A(n620), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n704) );
  AND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n703) );
  INV_X1 U735 ( .A(n703), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n661), .B(KEYINPUT81), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(KEYINPUT88), .ZN(n660) );
  INV_X1 U739 ( .A(KEYINPUT2), .ZN(n657) );
  OR2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  AND2_X1 U741 ( .A1(n403), .A2(KEYINPUT2), .ZN(n662) );
  INV_X1 U742 ( .A(n784), .ZN(n746) );
  NAND2_X1 U743 ( .A1(n662), .A2(n746), .ZN(n743) );
  NAND2_X1 U744 ( .A1(n757), .A2(G472), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(n478), .ZN(n667) );
  NOR2_X1 U746 ( .A1(n786), .A2(G952), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n446), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U750 ( .A(G104), .B(n671), .Z(G6) );
  NAND2_X1 U751 ( .A1(n690), .A2(n411), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(G146), .ZN(G48) );
  XNOR2_X1 U753 ( .A(G125), .B(KEYINPUT37), .ZN(n673) );
  XNOR2_X1 U754 ( .A(n674), .B(n673), .ZN(G27) );
  XNOR2_X1 U755 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n757), .A2(G469), .ZN(n680) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n681), .B(n682), .ZN(n683) );
  XOR2_X1 U760 ( .A(n684), .B(G101), .Z(G3) );
  AND2_X1 U761 ( .A1(n686), .A2(n685), .ZN(n688) );
  XNOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n687) );
  XNOR2_X1 U763 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U764 ( .A(G107), .B(n689), .ZN(G9) );
  XOR2_X1 U765 ( .A(G110), .B(n571), .Z(G12) );
  INV_X1 U766 ( .A(n690), .ZN(n691) );
  NOR2_X1 U767 ( .A1(n691), .A2(n369), .ZN(n695) );
  XOR2_X1 U768 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n693) );
  XNOR2_X1 U769 ( .A(n407), .B(KEYINPUT113), .ZN(n692) );
  XNOR2_X1 U770 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U771 ( .A(n695), .B(n694), .ZN(G30) );
  XOR2_X1 U772 ( .A(G143), .B(n696), .Z(G45) );
  NAND2_X1 U773 ( .A1(n698), .A2(n411), .ZN(n699) );
  XNOR2_X1 U774 ( .A(n699), .B(KEYINPUT114), .ZN(n700) );
  XNOR2_X1 U775 ( .A(G113), .B(n700), .ZN(G15) );
  NOR2_X1 U776 ( .A1(n701), .A2(n369), .ZN(n702) );
  XOR2_X1 U777 ( .A(G116), .B(n702), .Z(G18) );
  XOR2_X1 U778 ( .A(G134), .B(n703), .Z(G36) );
  XNOR2_X1 U779 ( .A(G140), .B(n704), .ZN(G42) );
  NOR2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n705) );
  XOR2_X1 U781 ( .A(KEYINPUT117), .B(n705), .Z(n709) );
  NAND2_X1 U782 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n716) );
  AND2_X1 U784 ( .A1(n711), .A2(n710), .ZN(n713) );
  AND2_X1 U785 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U786 ( .A(n714), .B(KEYINPUT118), .ZN(n715) );
  NOR2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U788 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n722) );
  INV_X1 U789 ( .A(n718), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U791 ( .A(n722), .B(n721), .ZN(n730) );
  NAND2_X1 U792 ( .A1(n724), .A2(n440), .ZN(n725) );
  XNOR2_X1 U793 ( .A(n725), .B(KEYINPUT115), .ZN(n726) );
  XNOR2_X1 U794 ( .A(KEYINPUT49), .B(n726), .ZN(n728) );
  NAND2_X1 U795 ( .A1(n728), .A2(n456), .ZN(n729) );
  OR2_X1 U796 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U797 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U798 ( .A(KEYINPUT51), .B(n733), .ZN(n734) );
  NOR2_X1 U799 ( .A1(n734), .A2(n740), .ZN(n735) );
  NOR2_X1 U800 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U801 ( .A(n737), .B(KEYINPUT52), .ZN(n738) );
  NOR2_X1 U802 ( .A1(n739), .A2(n738), .ZN(n741) );
  NOR2_X1 U803 ( .A1(n741), .A2(n359), .ZN(n751) );
  NOR2_X1 U804 ( .A1(n403), .A2(KEYINPUT2), .ZN(n742) );
  XNOR2_X1 U805 ( .A(n742), .B(KEYINPUT86), .ZN(n745) );
  INV_X1 U806 ( .A(n743), .ZN(n744) );
  NOR2_X1 U807 ( .A1(n745), .A2(n744), .ZN(n749) );
  XNOR2_X1 U808 ( .A(n747), .B(KEYINPUT87), .ZN(n748) );
  NAND2_X1 U809 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U810 ( .A(KEYINPUT53), .B(n753), .ZN(G75) );
  NAND2_X1 U811 ( .A1(n410), .A2(G478), .ZN(n755) );
  XOR2_X1 U812 ( .A(n755), .B(n405), .Z(n756) );
  NOR2_X1 U813 ( .A1(n761), .A2(n756), .ZN(G63) );
  NAND2_X1 U814 ( .A1(n410), .A2(G217), .ZN(n760) );
  XNOR2_X1 U815 ( .A(n758), .B(KEYINPUT122), .ZN(n759) );
  XNOR2_X1 U816 ( .A(n760), .B(n759), .ZN(n762) );
  NOR2_X1 U817 ( .A1(n762), .A2(n761), .ZN(G66) );
  XOR2_X1 U818 ( .A(KEYINPUT123), .B(n763), .Z(n766) );
  XNOR2_X1 U819 ( .A(G101), .B(n764), .ZN(n765) );
  XNOR2_X1 U820 ( .A(n766), .B(n765), .ZN(n768) );
  NOR2_X1 U821 ( .A1(n768), .A2(n767), .ZN(n777) );
  NAND2_X1 U822 ( .A1(n770), .A2(n403), .ZN(n774) );
  NAND2_X1 U823 ( .A1(G953), .A2(G224), .ZN(n771) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n771), .ZN(n772) );
  NAND2_X1 U825 ( .A1(n772), .A2(G898), .ZN(n773) );
  NAND2_X1 U826 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U827 ( .A(n775), .B(KEYINPUT124), .ZN(n776) );
  XNOR2_X1 U828 ( .A(n777), .B(n776), .ZN(G69) );
  XNOR2_X1 U829 ( .A(n778), .B(KEYINPUT125), .ZN(n779) );
  XNOR2_X1 U830 ( .A(n780), .B(n779), .ZN(n785) );
  XOR2_X1 U831 ( .A(G227), .B(n785), .Z(n781) );
  NAND2_X1 U832 ( .A1(n781), .A2(G900), .ZN(n782) );
  XNOR2_X1 U833 ( .A(KEYINPUT126), .B(n782), .ZN(n783) );
  NAND2_X1 U834 ( .A1(n783), .A2(G953), .ZN(n789) );
  XOR2_X1 U835 ( .A(n785), .B(n784), .Z(n787) );
  NAND2_X1 U836 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U837 ( .A1(n789), .A2(n788), .ZN(G72) );
  XOR2_X1 U838 ( .A(n406), .B(G122), .Z(G24) );
  XNOR2_X1 U839 ( .A(G131), .B(KEYINPUT127), .ZN(n792) );
  XNOR2_X1 U840 ( .A(n792), .B(n791), .ZN(G33) );
  XOR2_X1 U841 ( .A(G137), .B(n793), .Z(G39) );
endmodule

