//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(new_n206), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  NOR3_X1   g0017(.A1(new_n217), .A2(new_n213), .A3(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n215), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G226), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n210), .B2(new_n228), .C1(new_n203), .C2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n226), .B(new_n230), .C1(G97), .C2(G257), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(G1), .B2(G20), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n220), .B(new_n234), .C1(new_n216), .C2(new_n219), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT67), .B(G238), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n238), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n212), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n254), .B1(new_n217), .B2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n258), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n263), .A2(new_n213), .A3(G1), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n253), .A2(new_n212), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n272), .A2(new_n213), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT7), .ZN(new_n276));
  AOI211_X1 g0076(.A(new_n276), .B(G20), .C1(new_n269), .C2(new_n271), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n279), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT16), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n267), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n285), .A2(new_n286), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT75), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n269), .A2(new_n271), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n269), .B2(new_n271), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n213), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n287), .B1(new_n291), .B2(new_n276), .ZN(new_n292));
  OAI211_X1 g0092(.A(KEYINPUT16), .B(new_n281), .C1(new_n292), .C2(new_n203), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n266), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(G223), .A2(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n228), .A2(G1698), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n269), .A2(new_n295), .A3(new_n271), .A4(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT77), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n298), .B1(new_n297), .B2(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G1), .A3(G13), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(G232), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G274), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT78), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT78), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n304), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  INV_X1    g0118(.A(new_n314), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n306), .B2(new_n310), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n297), .A2(new_n299), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n318), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT18), .B1(new_n294), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n304), .B2(new_n315), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n321), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n284), .A2(new_n293), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(new_n265), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT17), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n265), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n317), .A2(new_n327), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n294), .A2(KEYINPUT17), .A3(new_n334), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n329), .A2(new_n338), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n346));
  INV_X1    g0146(.A(G150), .ZN(new_n347));
  INV_X1    g0147(.A(new_n280), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n213), .A2(G33), .ZN(new_n349));
  OAI221_X1 g0149(.A(new_n346), .B1(new_n347), .B2(new_n348), .C1(new_n261), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n254), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n264), .A2(new_n210), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n255), .A2(G50), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n350), .A2(new_n254), .B1(new_n210), .B2(new_n264), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT9), .B1(new_n357), .B2(new_n353), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G223), .A2(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G222), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n285), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n324), .C1(G77), .C2(new_n285), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n303), .A2(G226), .A3(new_n305), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n310), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n364), .A2(KEYINPUT68), .A3(new_n310), .A4(new_n365), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G200), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G190), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n359), .B(new_n374), .C1(KEYINPUT71), .C2(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n354), .A2(new_n355), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n357), .A2(KEYINPUT9), .A3(new_n353), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n371), .A3(new_n373), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n371), .A2(KEYINPUT71), .A3(new_n373), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n370), .A2(new_n318), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(new_n354), .C1(G179), .C2(new_n370), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n375), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AND4_X1   g0184(.A1(G226), .A2(new_n269), .A3(new_n271), .A4(new_n361), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n269), .A2(new_n271), .A3(G232), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n285), .A2(new_n388), .A3(G232), .A4(G1698), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n385), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n303), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n303), .A2(new_n305), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n310), .B1(new_n393), .B2(new_n229), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT13), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  INV_X1    g0196(.A(new_n394), .ZN(new_n397));
  INV_X1    g0197(.A(new_n391), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n398), .B(new_n385), .C1(new_n387), .C2(new_n389), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n396), .B(new_n397), .C1(new_n399), .C2(new_n303), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n400), .A3(G179), .ZN(new_n401));
  NAND2_X1  g0201(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT74), .A2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n395), .A2(new_n400), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n406), .B2(G169), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n318), .B(new_n404), .C1(new_n395), .C2(new_n400), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n203), .A2(G20), .ZN(new_n410));
  NOR3_X1   g0210(.A1(new_n410), .A2(G1), .A3(new_n263), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n255), .A2(G68), .B1(KEYINPUT12), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(KEYINPUT12), .B2(new_n411), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT73), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n410), .B1(new_n349), .B2(new_n222), .C1(new_n348), .C2(new_n210), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n254), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n418), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n406), .A2(G200), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n332), .C2(new_n406), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n263), .A2(G1), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G20), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G77), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n256), .A2(new_n222), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G20), .A2(G77), .ZN(new_n427));
  XOR2_X1   g0227(.A(KEYINPUT15), .B(G87), .Z(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n427), .B1(new_n348), .B2(new_n257), .C1(new_n429), .C2(new_n349), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n425), .B(new_n426), .C1(new_n254), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n361), .A2(G232), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n285), .B(new_n432), .C1(new_n229), .C2(new_n361), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(new_n324), .C1(G107), .C2(new_n285), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n310), .B1(new_n393), .B2(new_n223), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT70), .B(new_n310), .C1(new_n393), .C2(new_n223), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n431), .B(new_n440), .C1(new_n332), .C2(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(new_n431), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n439), .A2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n316), .B2(new_n439), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n422), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n345), .A2(new_n384), .A3(new_n419), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n424), .B2(G116), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n264), .A2(KEYINPUT83), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n267), .B(new_n424), .C1(G1), .C2(new_n268), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n253), .A2(new_n212), .B1(G20), .B2(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G283), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n457), .B(new_n213), .C1(G33), .C2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT20), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n456), .A2(KEYINPUT20), .A3(new_n459), .ZN(new_n461));
  OAI221_X1 g0261(.A(new_n454), .B1(new_n455), .B2(new_n452), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n324), .B1(new_n285), .B2(G303), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n361), .A2(G257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G264), .A2(G1698), .ZN(new_n467));
  AND4_X1   g0267(.A1(new_n269), .A2(new_n271), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n464), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G303), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n303), .B1(new_n272), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n285), .A2(new_n466), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(KEYINPUT82), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT79), .B1(new_n307), .B2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n307), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n308), .A2(G1), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n307), .A2(KEYINPUT5), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n478), .A2(G274), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n307), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n479), .B(new_n480), .C1(new_n482), .C2(new_n475), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G270), .A3(new_n303), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n474), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n463), .A2(new_n485), .A3(new_n316), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n462), .A3(G169), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT21), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n485), .A2(new_n462), .A3(new_n489), .A4(G169), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(G200), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n463), .C1(new_n332), .C2(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n225), .A2(new_n361), .ZN(new_n495));
  INV_X1    g0295(.A(G257), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(new_n495), .A3(new_n271), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n324), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n501), .A2(new_n481), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n483), .A2(G264), .A3(new_n303), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(G179), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n504), .A3(new_n481), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT85), .B1(new_n506), .B2(G169), .ZN(new_n507));
  AND4_X1   g0307(.A1(G179), .A2(new_n501), .A3(new_n504), .A4(new_n481), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n269), .A2(new_n271), .A3(new_n213), .A4(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT22), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT22), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n285), .A2(new_n514), .A3(new_n213), .A4(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(KEYINPUT84), .A2(KEYINPUT23), .A3(G107), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT84), .B1(new_n213), .B2(G107), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n213), .A2(new_n521), .B1(new_n522), .B2(new_n520), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n516), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT24), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n516), .A2(new_n526), .A3(new_n517), .A4(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n254), .ZN(new_n529));
  INV_X1    g0329(.A(new_n455), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(G107), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n423), .A2(G20), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g0333(.A(new_n533), .B(KEYINPUT25), .Z(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n505), .B(KEYINPUT86), .C1(new_n507), .C2(new_n508), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n511), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n528), .A2(new_n254), .B1(G107), .B2(new_n530), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n502), .A2(G190), .A3(new_n504), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n506), .A2(G200), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n534), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(G107), .B1(new_n275), .B2(new_n277), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n458), .A2(new_n532), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(KEYINPUT6), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n280), .A2(G77), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n543), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n254), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n424), .A2(G97), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n530), .A2(G97), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n481), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n269), .A2(new_n271), .A3(G244), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(G33), .B2(G283), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n559), .A2(G1698), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n285), .A2(G244), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n285), .B2(G250), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n560), .B(new_n562), .C1(new_n361), .C2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n557), .B1(new_n564), .B2(new_n324), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n483), .A2(new_n303), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G257), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n318), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n562), .A3(new_n457), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n285), .A2(G250), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n361), .B1(new_n571), .B2(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n324), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND4_X1   g0373(.A1(G179), .A2(new_n573), .A3(new_n567), .A4(new_n481), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n556), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n567), .A3(new_n481), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n553), .B1(new_n551), .B2(new_n254), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n573), .A2(new_n567), .A3(G190), .A4(new_n481), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n555), .A4(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT81), .ZN(new_n581));
  AND2_X1   g0381(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n582));
  NOR2_X1   g0382(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(G20), .B1(new_n584), .B2(new_n398), .ZN(new_n585));
  NOR3_X1   g0385(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n581), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n285), .A2(new_n213), .A3(G68), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n213), .B1(new_n589), .B2(new_n391), .ZN(new_n590));
  INV_X1    g0390(.A(new_n586), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(KEYINPUT81), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n458), .B2(new_n349), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n587), .A2(new_n588), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n254), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n428), .A2(new_n424), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n455), .A2(new_n429), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G274), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n479), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n225), .B1(new_n308), .B2(G1), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n303), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G238), .A2(G1698), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n223), .B2(G1698), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n285), .B1(G33), .B2(G116), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n607), .B2(new_n303), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n318), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G179), .B2(new_n608), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n600), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n330), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n332), .B(new_n604), .C1(new_n607), .C2(new_n303), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n455), .A2(new_n224), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n595), .A2(new_n615), .A3(new_n597), .A4(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n575), .A2(new_n580), .A3(new_n612), .A4(new_n618), .ZN(new_n619));
  NOR4_X1   g0419(.A1(new_n449), .A2(new_n494), .A3(new_n542), .A4(new_n619), .ZN(G372));
  AOI211_X1 g0420(.A(new_n596), .B(new_n616), .C1(new_n594), .C2(new_n254), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n615), .B1(new_n600), .B2(new_n611), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n541), .A2(new_n622), .A3(new_n575), .A4(new_n580), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n535), .A2(new_n509), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n491), .B2(new_n624), .ZN(new_n625));
  AOI211_X1 g0425(.A(new_n596), .B(new_n598), .C1(new_n594), .C2(new_n254), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n618), .B1(new_n626), .B2(new_n610), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT26), .B1(new_n627), .B2(new_n575), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n612), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n600), .A2(new_n611), .A3(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n576), .A2(G169), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n565), .A2(G179), .A3(new_n567), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n578), .B2(new_n555), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n612), .A4(new_n618), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n628), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n448), .B1(new_n625), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n383), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n329), .A2(new_n342), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n422), .A2(new_n442), .A3(new_n444), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n419), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n338), .A2(new_n343), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n375), .A2(new_n381), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G213), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT27), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n263), .A2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT88), .A3(new_n217), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n217), .A2(new_n213), .A3(G13), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(new_n656), .A3(new_n651), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT89), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n653), .A2(new_n656), .A3(new_n660), .A4(new_n651), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n650), .B(new_n657), .C1(new_n659), .C2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(KEYINPUT90), .B(G343), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n463), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n494), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n491), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n665), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n542), .ZN(new_n671));
  INV_X1    g0471(.A(new_n664), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n491), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n664), .B1(new_n538), .B2(new_n534), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n542), .A2(new_n675), .B1(new_n537), .B2(new_n664), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n624), .B1(new_n542), .B2(new_n491), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n664), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT91), .ZN(G399));
  INV_X1    g0483(.A(new_n218), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(G41), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n591), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n211), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n686), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n628), .A2(new_n632), .A3(new_n637), .ZN(new_n692));
  INV_X1    g0492(.A(new_n619), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n624), .A2(new_n491), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(new_n541), .A3(new_n694), .ZN(new_n695));
  AOI211_X1 g0495(.A(KEYINPUT29), .B(new_n672), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n638), .A2(KEYINPUT92), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n628), .A2(new_n632), .A3(new_n637), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n537), .A2(new_n491), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n537), .B2(new_n491), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n703), .A3(new_n623), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n664), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n696), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(new_n494), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n671), .A2(new_n707), .A3(new_n693), .A4(new_n664), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  AOI21_X1  g0509(.A(G179), .B1(new_n565), .B2(new_n567), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n485), .A3(new_n506), .A4(new_n608), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n565), .A2(new_n508), .A3(new_n567), .ZN(new_n713));
  INV_X1    g0513(.A(new_n608), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n474), .A3(new_n484), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n712), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n715), .ZN(new_n717));
  INV_X1    g0517(.A(new_n576), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n508), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n711), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n709), .B1(new_n720), .B2(new_n672), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n709), .A3(new_n672), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n708), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n706), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n691), .B1(new_n727), .B2(G1), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT94), .Z(G364));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT99), .Z(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n669), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n289), .ZN(new_n736));
  INV_X1    g0536(.A(new_n290), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n684), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(G45), .B2(new_n689), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT95), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n308), .B2(new_n248), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n285), .A2(new_n218), .A3(G355), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n743), .B(new_n744), .C1(G116), .C2(new_n218), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n212), .B1(G20), .B2(new_n318), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n732), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n652), .A2(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n686), .A2(G1), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n746), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n213), .A2(G179), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n330), .A2(G190), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n213), .A2(new_n316), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n332), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n272), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n332), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n213), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n757), .B(new_n763), .C1(G294), .C2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n332), .A2(new_n330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n758), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n758), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G311), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n758), .A2(new_n754), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n753), .A2(new_n772), .ZN(new_n778));
  INV_X1    g0578(.A(G329), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n768), .A2(new_n753), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n780), .B1(new_n783), .B2(G303), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n767), .A2(new_n771), .A3(new_n775), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n778), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n765), .A2(new_n458), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n769), .A2(new_n210), .B1(new_n773), .B2(new_n222), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n777), .A2(new_n203), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n285), .B1(new_n755), .B2(new_n532), .C1(new_n224), .C2(new_n781), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n202), .C2(new_n761), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n785), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n748), .B(new_n751), .C1(new_n752), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n735), .B1(KEYINPUT98), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(KEYINPUT98), .B2(new_n797), .ZN(new_n799));
  INV_X1    g0599(.A(new_n670), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n751), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(G330), .B2(new_n669), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  AOI21_X1  g0604(.A(new_n672), .B1(new_n692), .B2(new_n695), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n442), .A2(new_n672), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(new_n441), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT101), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n445), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(KEYINPUT101), .B1(new_n442), .B2(new_n444), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT102), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n445), .B2(new_n664), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n442), .A2(new_n444), .A3(new_n672), .A4(KEYINPUT102), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n805), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n726), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n750), .ZN(new_n819));
  INV_X1    g0619(.A(new_n777), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n760), .A2(G143), .B1(G150), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  INV_X1    g0622(.A(G159), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n821), .B1(new_n822), .B2(new_n769), .C1(new_n823), .C2(new_n773), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT34), .Z(new_n825));
  INV_X1    g0625(.A(new_n755), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G68), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n202), .B2(new_n765), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n739), .B1(new_n830), .B2(new_n778), .C1(new_n782), .C2(new_n210), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n755), .A2(new_n224), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n760), .B2(G294), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n778), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n835), .A2(new_n285), .A3(new_n789), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n836), .B1(new_n532), .B2(new_n782), .C1(new_n470), .C2(new_n769), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n452), .A2(new_n773), .B1(new_n777), .B2(new_n756), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT100), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n829), .A2(new_n831), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n746), .A2(new_n730), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n746), .B1(new_n222), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n811), .A2(new_n815), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n842), .B(new_n751), .C1(new_n731), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n819), .A2(new_n844), .ZN(G384));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n317), .A2(new_n327), .A3(new_n662), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n336), .B(new_n846), .C1(new_n294), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n327), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n326), .A2(new_n321), .A3(G179), .ZN(new_n852));
  INV_X1    g0652(.A(new_n662), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n339), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n855), .A2(KEYINPUT106), .A3(new_n846), .A4(new_n336), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n336), .B1(new_n294), .B2(new_n847), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT105), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n344), .A2(new_n339), .A3(new_n662), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n850), .A3(new_n856), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n281), .B1(new_n292), .B2(new_n203), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n283), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n293), .A2(new_n254), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n265), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n344), .A2(new_n662), .A3(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n870), .A2(new_n854), .B1(new_n294), .B2(new_n334), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n848), .B1(new_n872), .B2(new_n846), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n866), .A2(new_n874), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n542), .A2(new_n494), .A3(new_n619), .A4(new_n672), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n720), .A2(new_n709), .A3(new_n672), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n721), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n843), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n418), .A2(new_n672), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n409), .A2(new_n881), .A3(new_n418), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n409), .B2(new_n418), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n422), .B(new_n880), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n409), .A2(new_n418), .A3(new_n672), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT104), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n409), .A2(new_n888), .A3(new_n418), .A4(new_n672), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n879), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n875), .A2(new_n891), .A3(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n816), .B1(new_n708), .B2(new_n724), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n422), .A2(new_n880), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n419), .A2(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n882), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n887), .A2(new_n889), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT38), .B1(new_n871), .B2(new_n873), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n893), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n448), .A2(new_n725), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n904), .B(new_n905), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n883), .A2(new_n884), .A3(new_n672), .ZN(new_n908));
  INV_X1    g0708(.A(new_n901), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n874), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n900), .B1(new_n864), .B2(new_n865), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n908), .B(new_n910), .C1(new_n911), .C2(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n641), .A2(new_n853), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n890), .A2(new_n885), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n843), .B(new_n664), .C1(new_n625), .C2(new_n638), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n809), .A2(new_n672), .A3(new_n810), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n914), .B(new_n917), .C1(new_n900), .C2(new_n901), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n648), .B1(new_n706), .B2(new_n449), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n919), .B(new_n920), .Z(new_n921));
  XNOR2_X1  g0721(.A(new_n907), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n217), .B2(new_n652), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n452), .B1(new_n548), .B2(KEYINPUT35), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n924), .B(new_n214), .C1(KEYINPUT35), .C2(new_n548), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  OAI21_X1  g0726(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n689), .A2(new_n927), .B1(G50), .B2(new_n203), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n263), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n923), .A2(new_n926), .A3(new_n929), .ZN(G367));
  AND2_X1   g0730(.A1(new_n575), .A2(new_n580), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n672), .A2(new_n556), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(KEYINPUT108), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT109), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n575), .B2(new_n664), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n635), .A2(KEYINPUT109), .A3(new_n672), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n674), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(KEYINPUT42), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT42), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n935), .A2(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(new_n674), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n575), .B1(new_n946), .B2(new_n537), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n664), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n621), .A2(new_n664), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n630), .A2(new_n631), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n627), .B2(new_n952), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT107), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n948), .B(new_n950), .C1(KEYINPUT43), .C2(new_n955), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT110), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT110), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n957), .A2(new_n962), .A3(new_n959), .A4(new_n958), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n679), .A2(new_n946), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n749), .A2(G1), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT44), .B1(new_n942), .B2(new_n681), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n946), .A2(new_n971), .A3(new_n664), .A4(new_n680), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n942), .A2(new_n681), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n942), .B2(new_n681), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n970), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n670), .B(new_n677), .Z(new_n978));
  NAND3_X1  g0778(.A1(new_n727), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n979), .A2(new_n727), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n685), .B(KEYINPUT41), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n969), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n961), .A2(new_n965), .A3(new_n963), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n967), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n740), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n747), .B1(new_n218), .B2(new_n429), .C1(new_n986), .C2(new_n244), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G283), .A2(new_n774), .B1(new_n826), .B2(G97), .ZN(new_n988));
  INV_X1    g0788(.A(G294), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n989), .B2(new_n777), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n738), .B1(new_n532), .B2(new_n765), .C1(new_n991), .C2(new_n778), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(G303), .C2(new_n760), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT46), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n783), .B2(G116), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n993), .B1(new_n834), .B2(new_n769), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT111), .ZN(new_n998));
  INV_X1    g0798(.A(new_n781), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G143), .A2(new_n770), .B1(new_n999), .B2(G58), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n822), .B2(new_n778), .C1(new_n823), .C2(new_n777), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n285), .B1(new_n755), .B2(new_n222), .C1(new_n761), .C2(new_n347), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n773), .A2(new_n210), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n765), .A2(new_n203), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n751), .B(new_n987), .C1(new_n1007), .C2(new_n752), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT112), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n734), .B2(new_n954), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  OR2_X1    g0811(.A1(new_n727), .A2(new_n978), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n727), .A2(new_n978), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n685), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n978), .A2(new_n968), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n740), .B1(new_n241), .B2(new_n308), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n687), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n218), .A3(new_n285), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n257), .A2(G50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1017), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(G68), .A2(G77), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n308), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1019), .A2(new_n1024), .B1(new_n532), .B2(new_n684), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n747), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n751), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT113), .Z(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n774), .B1(new_n820), .B2(G311), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT115), .B(G322), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n769), .B2(new_n1030), .C1(new_n991), .C2(new_n761), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT48), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n756), .B2(new_n765), .C1(new_n989), .C2(new_n781), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n786), .A2(G326), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n739), .B1(G116), .B2(new_n826), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G68), .A2(new_n774), .B1(new_n786), .B2(G150), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n458), .B2(new_n755), .C1(new_n823), .C2(new_n769), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n261), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n820), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n429), .A2(new_n765), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G50), .B2(new_n760), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n999), .A2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1046), .A3(new_n739), .A4(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1039), .A2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1028), .B1(new_n676), .B2(new_n734), .C1(new_n1049), .C2(new_n752), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1014), .A2(new_n1015), .A3(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n977), .A2(new_n678), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n970), .A2(new_n972), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n679), .C1(new_n975), .C2(new_n976), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n1013), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n685), .A3(new_n979), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n1054), .A3(new_n968), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n747), .B1(new_n458), .B2(new_n218), .C1(new_n986), .C2(new_n251), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n760), .A2(G159), .B1(new_n770), .B2(G150), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n739), .B1(new_n257), .B2(new_n773), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G50), .A2(new_n820), .B1(new_n786), .B2(G143), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n766), .A2(G77), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n203), .C2(new_n781), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1061), .A2(new_n832), .A3(new_n1062), .A4(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT116), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G294), .A2(new_n774), .B1(new_n820), .B2(G303), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n756), .B2(new_n781), .C1(new_n778), .C2(new_n1030), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n285), .B(new_n1069), .C1(G116), .C2(new_n766), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n760), .A2(G311), .B1(new_n770), .B2(G317), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT52), .Z(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n532), .C2(new_n755), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n750), .B1(new_n1074), .B2(new_n746), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n732), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1059), .B(new_n1075), .C1(new_n942), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1058), .A2(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1057), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  OAI211_X1 g0880(.A(new_n894), .B(G330), .C1(new_n897), .C2(new_n898), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n908), .B1(new_n914), .B2(new_n917), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT39), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n859), .A2(new_n850), .A3(new_n856), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT105), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n850), .A2(new_n856), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT38), .B1(new_n1089), .B2(new_n862), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1090), .B2(new_n900), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1083), .B1(new_n1091), .B2(new_n910), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n908), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1090), .B2(new_n900), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n897), .A2(new_n898), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n664), .B(new_n843), .C1(new_n700), .C2(new_n704), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n916), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1082), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1083), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n910), .B1(new_n911), .B2(KEYINPUT39), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1096), .A2(new_n916), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1093), .B(new_n875), .C1(new_n1103), .C2(new_n1095), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(new_n1104), .A3(new_n1081), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n448), .A2(G330), .A3(new_n725), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n648), .C1(new_n706), .C2(new_n449), .ZN(new_n1107));
  INV_X1    g0907(.A(G330), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n885), .B(new_n890), .C1(new_n879), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1081), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n917), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1103), .A2(new_n1081), .A3(new_n1109), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1099), .A2(new_n1105), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT117), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1107), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1099), .A2(new_n1105), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n685), .B(new_n1114), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1101), .A2(new_n730), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n778), .A2(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n285), .B1(new_n755), .B2(new_n210), .C1(new_n822), .C2(new_n777), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G159), .C2(new_n766), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n761), .A2(new_n830), .B1(new_n773), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT53), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n781), .B2(new_n347), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n999), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G128), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1127), .B(new_n1134), .C1(new_n1135), .C2(new_n769), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT118), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n769), .A2(new_n756), .B1(new_n777), .B2(new_n532), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G97), .B2(new_n774), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT119), .Z(new_n1140));
  NAND2_X1  g0940(.A1(new_n760), .A2(G116), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n1064), .A3(new_n272), .A4(new_n827), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G87), .B2(new_n783), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1140), .B(new_n1143), .C1(new_n989), .C2(new_n778), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1137), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n750), .B1(new_n1145), .B2(new_n746), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1123), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n261), .B2(new_n841), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1121), .B2(new_n968), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1122), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G378));
  NAND3_X1  g0951(.A1(new_n892), .A2(new_n903), .A3(G330), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT55), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n384), .B(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n853), .B1(new_n357), .B2(new_n353), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT56), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1154), .B(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1156), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1154), .B(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1160), .A2(new_n892), .A3(G330), .A4(new_n903), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n919), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n919), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1163), .A2(new_n1165), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n686), .B1(new_n1166), .B2(KEYINPUT57), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1158), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1168), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1157), .A2(new_n730), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n841), .A2(new_n210), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G58), .A2(new_n826), .B1(new_n786), .B2(G283), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n458), .B2(new_n777), .C1(new_n429), .C2(new_n773), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1004), .B(new_n1179), .C1(G116), .C2(new_n770), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n738), .A2(new_n307), .A3(new_n1047), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT120), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(new_n532), .C2(new_n761), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT58), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n765), .A2(new_n347), .B1(new_n769), .B2(new_n1124), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n760), .A2(G128), .B1(new_n999), .B2(new_n1128), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n822), .B2(new_n773), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G132), .C2(new_n820), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT59), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G41), .B1(new_n786), .B2(G124), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G33), .B1(new_n826), .B2(G159), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G41), .B1(new_n739), .B2(G33), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1184), .B(new_n1192), .C1(G50), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n750), .B1(new_n1194), .B2(new_n746), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1176), .A2(new_n1177), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n968), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1175), .A2(new_n1199), .ZN(G375));
  AOI21_X1  g1000(.A(new_n969), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT122), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n777), .A2(new_n452), .B1(new_n778), .B2(new_n470), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n783), .B2(G97), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n774), .A2(G107), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n272), .B1(new_n755), .B2(new_n222), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1206), .B(new_n1044), .C1(G283), .C2(new_n760), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G294), .B2(new_n770), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n760), .A2(G137), .B1(G150), .B2(new_n774), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n1135), .B2(new_n778), .C1(new_n782), .C2(new_n823), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1129), .A2(new_n777), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n739), .B1(new_n830), .B2(new_n769), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n765), .A2(new_n210), .B1(new_n202), .B2(new_n755), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n746), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n841), .A2(new_n203), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n751), .A3(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT121), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1095), .B2(new_n730), .ZN(new_n1220));
  OR3_X1    g1020(.A1(new_n1201), .A2(new_n1202), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1202), .B1(new_n1201), .B2(new_n1220), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1111), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1225), .B2(new_n982), .ZN(G381));
  NAND3_X1  g1026(.A1(new_n1175), .A2(new_n1150), .A3(new_n1199), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(G396), .A3(G393), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n985), .A2(new_n1079), .A3(new_n1010), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(G384), .A3(G381), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(G407));
  OAI211_X1 g1031(.A(G407), .B(G213), .C1(new_n663), .C2(new_n1227), .ZN(G409));
  XNOR2_X1  g1032(.A(G393), .B(new_n803), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n985), .A2(new_n1079), .A3(new_n1010), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1079), .B1(new_n985), .B2(new_n1010), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G387), .A2(G390), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1233), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1229), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n663), .A2(new_n650), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1166), .A2(new_n981), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1243), .A2(new_n1199), .A3(new_n1149), .A4(new_n1122), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1196), .B1(new_n1173), .B2(new_n969), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1242), .B(new_n1244), .C1(new_n1246), .C2(new_n1150), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1113), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1224), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1111), .A2(new_n1107), .A3(new_n1112), .A4(KEYINPUT60), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1250), .A3(new_n685), .A4(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1223), .A2(G384), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(G384), .B1(new_n1223), .B2(new_n1252), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT123), .B1(new_n1247), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1244), .A2(new_n1242), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT123), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .A4(new_n1256), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT62), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1241), .A2(G2897), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT125), .Z(new_n1266));
  NAND2_X1  g1066(.A1(new_n1256), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1266), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1150), .B1(new_n1175), .B2(new_n1199), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1267), .B(new_n1269), .C1(new_n1270), .C2(new_n1260), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1270), .A2(new_n1260), .A3(new_n1257), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1271), .B(new_n1272), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1240), .B1(new_n1264), .B2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(KEYINPUT124), .B(KEYINPUT63), .Z(new_n1277));
  NAND3_X1  g1077(.A1(new_n1258), .A2(new_n1263), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1240), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(KEYINPUT63), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(G405));
  NOR2_X1   g1083(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1236), .A2(new_n1239), .A3(KEYINPUT127), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1240), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1284), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1236), .A2(new_n1239), .A3(KEYINPUT127), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1259), .A2(new_n1293), .A3(new_n1227), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1287), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1287), .B2(new_n1292), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


