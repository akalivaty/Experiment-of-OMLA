//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G162gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n207), .A2(new_n208), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(KEYINPUT77), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G155gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n208), .B1(new_n218), .B2(G162gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n205), .A2(new_n210), .A3(new_n212), .A4(new_n206), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n219), .A2(KEYINPUT78), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT77), .B(G155gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT2), .B1(new_n223), .B2(new_n209), .ZN(new_n224));
  AND4_X1   g023(.A1(new_n210), .A2(new_n205), .A3(new_n212), .A4(new_n206), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n214), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  XOR2_X1   g027(.A(G113gat), .B(G120gat), .Z(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G113gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n236), .A3(G120gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n233), .A2(G120gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n230), .A3(new_n228), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT69), .B(G113gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n243), .B2(G120gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(new_n238), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n232), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n202), .B1(new_n227), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT78), .B1(new_n219), .B2(new_n220), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n225), .A3(new_n222), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n213), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n230), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n244), .B2(new_n238), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n240), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT70), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n231), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT4), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n246), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  AOI211_X1 g057(.A(KEYINPUT3), .B(new_n213), .C1(new_n248), .C2(new_n249), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n247), .B(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n227), .A2(new_n246), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n250), .A2(new_n255), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI22_X1  g065(.A1(new_n260), .A2(new_n262), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT0), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G85gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n247), .A2(new_n256), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n257), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n274), .A3(new_n246), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(KEYINPUT5), .A3(new_n261), .A4(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n267), .A2(new_n276), .ZN(new_n281));
  INV_X1    g080(.A(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n271), .B(KEYINPUT81), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n276), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT26), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n290), .A2(new_n295), .A3(new_n291), .A4(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(G169gat), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n291), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n288), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT27), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT27), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n307), .B1(new_n312), .B2(new_n308), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n302), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n316), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT23), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n288), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n316), .A2(G169gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G176gat), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT66), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n297), .A2(new_n298), .B1(new_n318), .B2(KEYINPUT23), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n300), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT64), .B(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n321), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G183gat), .B(G190gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n334), .B(new_n336), .C1(new_n337), .C2(new_n335), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n303), .A2(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n308), .A2(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT24), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n290), .A2(KEYINPUT23), .A3(new_n292), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n344), .A3(new_n336), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT25), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n315), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(KEYINPUT75), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n351), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G197gat), .B(G204gat), .ZN(new_n359));
  INV_X1    g158(.A(G211gat), .ZN(new_n360));
  INV_X1    g159(.A(G218gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(KEYINPUT22), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G211gat), .B(G218gat), .Z(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n365), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT74), .B1(new_n348), .B2(new_n353), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  AOI211_X1 g168(.A(KEYINPUT74), .B(new_n353), .C1(new_n348), .C2(new_n349), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n366), .A2(new_n371), .A3(new_n377), .A4(new_n374), .ZN(new_n378));
  AND4_X1   g177(.A1(new_n280), .A2(new_n287), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n374), .B1(new_n366), .B2(new_n371), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT37), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n366), .B2(new_n371), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n380), .B(KEYINPUT38), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n374), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n350), .A2(new_n351), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n354), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n357), .A2(new_n389), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n365), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT75), .B1(new_n348), .B2(new_n353), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n317), .A2(new_n319), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(new_n300), .B1(new_n331), .B2(new_n321), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n338), .B1(new_n396), .B2(new_n330), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(new_n326), .B1(KEYINPUT25), .B2(new_n346), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n398), .B2(new_n315), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n399), .B2(new_n353), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n367), .B1(new_n400), .B2(new_n352), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n387), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n383), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n366), .A2(new_n371), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n402), .A2(new_n403), .B1(new_n404), .B2(KEYINPUT37), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT38), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT83), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n358), .A2(new_n367), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT37), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n406), .B(new_n410), .C1(new_n381), .C2(new_n383), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n379), .A2(new_n386), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n365), .B1(new_n274), .B2(new_n349), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT3), .B1(new_n365), .B2(new_n349), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n250), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT79), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n414), .B2(new_n250), .ZN(new_n418));
  AND2_X1   g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n419), .C1(new_n413), .C2(new_n415), .ZN(new_n422));
  AOI21_X1  g221(.A(G22gat), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(G22gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT31), .B(G50gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n429), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n424), .A2(new_n430), .A3(new_n425), .A4(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n260), .A2(new_n262), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n264), .A2(new_n265), .A3(new_n261), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(KEYINPUT39), .A3(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT82), .B(KEYINPUT39), .Z(new_n438));
  NAND3_X1  g237(.A1(new_n260), .A2(new_n262), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n284), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n286), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n441), .B2(new_n440), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n376), .A2(new_n444), .A3(new_n378), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT30), .A4(new_n374), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n402), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n434), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n412), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT6), .B1(new_n281), .B2(new_n282), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n277), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n280), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n445), .A3(new_n447), .ZN(new_n454));
  NAND2_X1  g253(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n398), .A2(new_n246), .A3(new_n315), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n348), .A2(new_n255), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n460), .A3(G227gat), .A4(G233gat), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n458), .B1(new_n461), .B2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(new_n461), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(KEYINPUT33), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n458), .A2(KEYINPUT71), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(KEYINPUT71), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(KEYINPUT33), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n459), .A2(new_n460), .ZN(new_n469));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470));
  AND2_X1   g269(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n464), .A2(new_n468), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n464), .B2(new_n468), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n455), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n468), .ZN(new_n480));
  INV_X1    g279(.A(new_n475), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n483));
  INV_X1    g282(.A(new_n455), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n476), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n454), .A2(new_n434), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n432), .A2(new_n482), .A3(new_n433), .A4(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n454), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n448), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n432), .A2(new_n433), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n477), .A2(new_n478), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT35), .B1(new_n287), .B2(new_n280), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n450), .A2(new_n486), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(KEYINPUT13), .Z(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  AND2_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G29gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n505));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI221_X1 g316(.A(new_n513), .B1(new_n514), .B2(new_n510), .C1(G1gat), .C2(new_n511), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n520), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n509), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n523), .ZN(new_n525));
  INV_X1    g324(.A(new_n509), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n496), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n519), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n509), .A2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n507), .B2(new_n508), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n522), .A2(new_n509), .A3(new_n523), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT18), .A4(new_n495), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n495), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT86), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT12), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n536), .B(new_n539), .C1(new_n540), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n540), .A3(new_n535), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(new_n539), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n535), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n546), .A2(KEYINPUT87), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT87), .B1(new_n546), .B2(new_n551), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n494), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n557), .A2(G85gat), .A3(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G99gat), .B(G106gat), .ZN(new_n560));
  XOR2_X1   g359(.A(KEYINPUT97), .B(G85gat), .Z(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT98), .B(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n561), .A2(new_n562), .B1(KEYINPUT8), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n559), .A2(new_n564), .ZN(new_n567));
  INV_X1    g366(.A(new_n560), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(KEYINPUT99), .A3(new_n565), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n566), .B(new_n570), .C1(new_n530), .C2(new_n532), .ZN(new_n571));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT93), .Z(new_n573));
  INV_X1    g372(.A(KEYINPUT41), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n566), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n509), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n571), .A2(new_n577), .A3(new_n308), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n308), .B1(new_n571), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n361), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n571), .A2(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G190gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(new_n577), .A3(new_n308), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(G218gat), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n573), .A2(new_n574), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  NAND4_X1  g389(.A1(new_n580), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G64gat), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n598), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT88), .B1(new_n604), .B2(new_n602), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(KEYINPUT88), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n602), .B1(new_n604), .B2(new_n601), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT89), .B1(new_n597), .B2(G64gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n598), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n600), .A2(KEYINPUT89), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n608), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G231gat), .ZN(new_n620));
  INV_X1    g419(.A(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n617), .B(new_n618), .C1(new_n620), .C2(new_n621), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n623), .B2(new_n624), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n596), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(new_n596), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n626), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n595), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n525), .A2(new_n521), .B1(new_n618), .B2(new_n617), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n632), .A3(new_n595), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n637), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n633), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n590), .B1(new_n589), .B2(new_n591), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n593), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n615), .A2(new_n616), .ZN(new_n647));
  AOI22_X1  g446(.A1(new_n570), .A2(new_n566), .B1(new_n647), .B2(new_n608), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n617), .B1(new_n565), .B2(new_n569), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n576), .A2(KEYINPUT10), .A3(new_n608), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n648), .A2(new_n653), .A3(new_n649), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n656), .B(new_n657), .Z(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT100), .B1(new_n652), .B2(new_n653), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  INV_X1    g461(.A(new_n653), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n662), .B(new_n663), .C1(new_n650), .C2(new_n651), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n655), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n658), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n555), .A2(new_n645), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n453), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT101), .B(G1gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1324gat));
  NAND2_X1  g470(.A1(new_n589), .A2(new_n591), .ZN(new_n672));
  INV_X1    g471(.A(new_n590), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n639), .A2(new_n642), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n592), .A4(new_n667), .ZN(new_n676));
  NOR4_X1   g475(.A1(new_n494), .A2(new_n489), .A3(new_n554), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT103), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT102), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n682), .B(new_n684), .C1(new_n510), .C2(new_n677), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n485), .A2(new_n479), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n668), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n491), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n668), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n668), .A2(new_n490), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n592), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n665), .A2(new_n666), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n659), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n675), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g496(.A1(new_n555), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n279), .B1(new_n451), .B2(new_n277), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n501), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n593), .A2(new_n644), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n494), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n434), .B1(new_n448), .B2(new_n699), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n686), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n412), .B2(new_n449), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n493), .A2(new_n488), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n694), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n546), .A2(new_n551), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n697), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n453), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n701), .A2(new_n713), .ZN(G1328gat));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n497), .A3(new_n448), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT46), .Z(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n489), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  OAI21_X1  g517(.A(G43gat), .B1(new_n712), .B2(new_n686), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n720), .A3(new_n491), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g522(.A(G50gat), .B1(new_n712), .B2(new_n490), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n698), .A2(new_n725), .A3(new_n434), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g527(.A1(new_n450), .A2(new_n486), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n493), .A2(new_n488), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n711), .ZN(new_n732));
  AND4_X1   g531(.A1(new_n731), .A2(new_n732), .A3(new_n645), .A4(new_n696), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n699), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n448), .B1(new_n736), .B2(new_n599), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n599), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  INV_X1    g540(.A(new_n686), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n688), .A2(G71gat), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n743), .A2(G71gat), .B1(new_n733), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n733), .A2(new_n434), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT106), .B(G78gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n703), .B1(new_n729), .B2(new_n730), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n675), .A2(new_n711), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  INV_X1    g554(.A(new_n753), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n494), .A2(new_n755), .A3(new_n703), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT108), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n731), .A2(new_n694), .A3(new_n753), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n755), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n751), .B1(new_n758), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n752), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n761), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n754), .A2(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n561), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n453), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n763), .A2(new_n696), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n756), .A2(new_n667), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n704), .A2(new_n709), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n704), .A2(new_n709), .A3(KEYINPUT107), .A4(new_n771), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n699), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n768), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n770), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n770), .A2(KEYINPUT110), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1336gat));
  NOR3_X1   g581(.A1(new_n489), .A2(new_n667), .A3(G92gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT112), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n710), .A2(new_n448), .A3(new_n771), .ZN(new_n786));
  INV_X1    g585(.A(new_n562), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n448), .A3(new_n775), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(new_n783), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n760), .B2(new_n764), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT111), .B1(new_n795), .B2(KEYINPUT52), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n790), .B2(new_n787), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n789), .B1(new_n796), .B2(new_n800), .ZN(G1337gat));
  NOR2_X1   g600(.A1(new_n688), .A2(G99gat), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n763), .A2(new_n696), .A3(new_n767), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n774), .A2(new_n742), .A3(new_n775), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G99gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n490), .A2(new_n667), .A3(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n765), .A2(new_n766), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI21_X1  g608(.A(G106gat), .B1(new_n772), .B2(new_n490), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n774), .A2(new_n434), .A3(new_n775), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n760), .A2(new_n764), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n812), .A2(G106gat), .B1(new_n813), .B2(new_n807), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n814), .B2(new_n809), .ZN(G1339gat));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n645), .A2(new_n816), .A3(new_n732), .A4(new_n667), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n676), .B2(new_n711), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n661), .A2(new_n664), .A3(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n650), .A2(new_n663), .A3(new_n651), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n666), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n661), .ZN(new_n826));
  INV_X1    g625(.A(new_n664), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n652), .B2(new_n653), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n658), .B1(new_n830), .B2(new_n822), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n825), .A2(new_n832), .A3(new_n711), .A4(new_n659), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n526), .B1(new_n525), .B2(new_n521), .ZN(new_n834));
  INV_X1    g633(.A(new_n496), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n534), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n533), .A2(new_n534), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(G229gat), .A3(G233gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n834), .A2(new_n534), .A3(KEYINPUT114), .A4(new_n835), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(KEYINPUT115), .A3(new_n544), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n536), .A2(new_n539), .A3(new_n545), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n842), .B2(new_n544), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n696), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n703), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n825), .A2(new_n832), .A3(new_n659), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n694), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n675), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n819), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n453), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n487), .A2(new_n448), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n243), .A3(new_n711), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n490), .B1(new_n819), .B2(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT116), .B(new_n490), .C1(new_n819), .C2(new_n854), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n448), .A2(new_n453), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n688), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n865), .B2(new_n869), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n554), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n860), .B1(new_n872), .B2(new_n233), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n859), .B2(new_n696), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n870), .A2(new_n871), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n696), .A2(G120gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G1341gat));
  INV_X1    g676(.A(G127gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n878), .A3(new_n675), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n870), .A2(new_n871), .A3(new_n643), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n878), .ZN(G1342gat));
  INV_X1    g680(.A(G134gat), .ZN(new_n882));
  AND4_X1   g681(.A1(new_n882), .A2(new_n856), .A3(new_n857), .A4(new_n694), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT56), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n870), .A2(new_n871), .A3(new_n703), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n882), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n434), .C1(new_n819), .C2(new_n854), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n868), .A2(new_n742), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n842), .A2(new_n544), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n843), .A3(new_n844), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT118), .B1(new_n895), .B2(new_n667), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n847), .A2(new_n696), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n898), .C1(new_n554), .C2(new_n851), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n703), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n703), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n853), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n643), .ZN(new_n905));
  INV_X1    g704(.A(new_n819), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n490), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n711), .B(new_n891), .C1(new_n907), .C2(new_n887), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n686), .A2(KEYINPUT121), .A3(new_n434), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT121), .B1(new_n686), .B2(new_n434), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n489), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n819), .A2(new_n854), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(KEYINPUT120), .A3(new_n699), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n855), .B2(new_n453), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n554), .A2(G141gat), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n908), .A2(G141gat), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n703), .A2(new_n895), .A3(new_n851), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n900), .B2(new_n901), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n675), .B1(new_n921), .B2(new_n903), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n434), .B1(new_n922), .B2(new_n819), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n890), .B1(new_n923), .B2(KEYINPUT57), .ZN(new_n924));
  INV_X1    g723(.A(new_n554), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n203), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n916), .A2(new_n917), .ZN(new_n927));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n918), .A2(new_n919), .B1(new_n926), .B2(new_n929), .ZN(G1344gat));
  OAI211_X1 g729(.A(new_n696), .B(new_n891), .C1(new_n907), .C2(new_n887), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n204), .A2(KEYINPUT59), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n434), .B1(new_n819), .B2(new_n854), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(KEYINPUT57), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n675), .B1(new_n900), .B2(new_n853), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n676), .A2(new_n925), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n887), .B(new_n434), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n868), .A2(new_n742), .A3(new_n667), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G148gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT123), .B1(new_n941), .B2(KEYINPUT59), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n943), .B(new_n944), .C1(new_n940), .C2(G148gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n933), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n916), .A2(new_n204), .A3(new_n696), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1345gat));
  NAND3_X1  g747(.A1(new_n916), .A2(new_n223), .A3(new_n675), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n924), .A2(new_n675), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n223), .ZN(G1346gat));
  AOI21_X1  g750(.A(G162gat), .B1(new_n916), .B2(new_n694), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n703), .A2(new_n209), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n924), .B2(new_n953), .ZN(G1347gat));
  NAND2_X1  g753(.A1(new_n448), .A2(new_n453), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n855), .A2(new_n487), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n711), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n688), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n959), .B1(new_n863), .B2(new_n864), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n554), .A2(new_n297), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(G1348gat));
  AOI21_X1  g761(.A(G176gat), .B1(new_n956), .B2(new_n696), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n667), .A2(new_n331), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n960), .B2(new_n964), .ZN(G1349gat));
  AOI21_X1  g764(.A(new_n303), .B1(new_n960), .B2(new_n675), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n955), .A2(new_n487), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n675), .A2(new_n312), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n967), .B(new_n968), .C1(new_n819), .C2(new_n854), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(KEYINPUT125), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n966), .A2(new_n971), .A3(KEYINPUT60), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT60), .B1(new_n966), .B2(new_n971), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1350gat));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  AOI211_X1 g774(.A(new_n703), .B(new_n959), .C1(new_n863), .C2(new_n864), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n976), .B2(new_n308), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n865), .A2(new_n694), .A3(new_n958), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n975), .B(new_n981), .C1(new_n976), .C2(new_n308), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n956), .A2(new_n308), .A3(new_n694), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(G1351gat));
  INV_X1    g783(.A(new_n934), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n742), .A2(new_n955), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n711), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n935), .A2(new_n938), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n986), .B(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n925), .A2(G197gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(G1352gat));
  OAI21_X1  g794(.A(G204gat), .B1(new_n992), .B2(new_n667), .ZN(new_n996));
  OR2_X1    g795(.A1(new_n667), .A2(G204gat), .ZN(new_n997));
  OAI21_X1  g796(.A(KEYINPUT62), .B1(new_n987), .B2(new_n997), .ZN(new_n998));
  OR3_X1    g797(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n988), .A2(new_n360), .A3(new_n675), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n990), .A2(new_n675), .A3(new_n991), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  OAI21_X1  g804(.A(G218gat), .B1(new_n992), .B2(new_n703), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n361), .A3(new_n694), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1355gat));
endmodule


