

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781;

  AND2_X1 U384 ( .A1(n393), .A2(n414), .ZN(n411) );
  BUF_X1 U385 ( .A(n720), .Z(n364) );
  NAND2_X1 U386 ( .A1(n441), .A2(n439), .ZN(n362) );
  BUF_X1 U387 ( .A(n687), .Z(n365) );
  XNOR2_X1 U388 ( .A(n452), .B(n451), .ZN(n720) );
  NAND2_X1 U389 ( .A1(n568), .A2(n623), .ZN(n452) );
  XNOR2_X1 U390 ( .A(n603), .B(KEYINPUT1), .ZN(n687) );
  BUF_X1 U391 ( .A(n557), .Z(n693) );
  XNOR2_X1 U392 ( .A(n453), .B(G469), .ZN(n603) );
  OR2_X1 U393 ( .A1(n738), .A2(G902), .ZN(n453) );
  XNOR2_X1 U394 ( .A(n766), .B(n490), .ZN(n526) );
  XNOR2_X1 U395 ( .A(n496), .B(G140), .ZN(n497) );
  XNOR2_X1 U396 ( .A(G116), .B(G113), .ZN(n460) );
  INV_X2 U397 ( .A(G953), .ZN(n769) );
  NOR2_X1 U398 ( .A1(n363), .A2(n362), .ZN(n438) );
  AND2_X2 U399 ( .A1(n577), .A2(KEYINPUT34), .ZN(n363) );
  OR2_X2 U400 ( .A1(n657), .A2(G902), .ZN(n527) );
  XNOR2_X1 U401 ( .A(G143), .B(G113), .ZN(n533) );
  XNOR2_X1 U402 ( .A(n461), .B(n460), .ZN(n520) );
  INV_X1 U403 ( .A(n680), .ZN(n678) );
  XNOR2_X1 U404 ( .A(n563), .B(n562), .ZN(n661) );
  XNOR2_X2 U405 ( .A(n403), .B(n385), .ZN(n369) );
  NAND2_X2 U406 ( .A1(n413), .A2(n412), .ZN(n742) );
  NAND2_X2 U407 ( .A1(n411), .A2(n430), .ZN(n413) );
  NAND2_X2 U408 ( .A1(n415), .A2(n372), .ZN(n412) );
  INV_X2 U409 ( .A(KEYINPUT3), .ZN(n459) );
  INV_X2 U410 ( .A(G125), .ZN(n454) );
  NAND2_X2 U411 ( .A1(n409), .A2(n407), .ZN(n587) );
  XNOR2_X2 U412 ( .A(n550), .B(KEYINPUT4), .ZN(n489) );
  XNOR2_X2 U413 ( .A(n424), .B(n489), .ZN(n766) );
  NOR2_X1 U414 ( .A1(n597), .A2(n519), .ZN(n688) );
  INV_X1 U415 ( .A(KEYINPUT48), .ZN(n446) );
  XNOR2_X1 U416 ( .A(G104), .B(G110), .ZN(n463) );
  XNOR2_X1 U417 ( .A(n643), .B(KEYINPUT46), .ZN(n448) );
  AND2_X1 U418 ( .A1(n661), .A2(n408), .ZN(n407) );
  INV_X1 U419 ( .A(n673), .ZN(n366) );
  AND2_X1 U420 ( .A1(n604), .A2(n603), .ZN(n456) );
  AND2_X1 U421 ( .A1(n687), .A2(n688), .ZN(n568) );
  XNOR2_X1 U422 ( .A(n527), .B(G472), .ZN(n557) );
  XNOR2_X1 U423 ( .A(n459), .B(G119), .ZN(n461) );
  XNOR2_X1 U424 ( .A(n463), .B(G107), .ZN(n752) );
  INV_X2 U425 ( .A(KEYINPUT70), .ZN(n488) );
  NAND2_X1 U426 ( .A1(n413), .A2(n412), .ZN(n367) );
  BUF_X1 U427 ( .A(n755), .Z(n368) );
  XNOR2_X1 U428 ( .A(n520), .B(n462), .ZN(n755) );
  BUF_X1 U429 ( .A(n664), .Z(n370) );
  BUF_X1 U430 ( .A(n781), .Z(n371) );
  XNOR2_X2 U431 ( .A(n625), .B(n387), .ZN(n455) );
  XNOR2_X1 U432 ( .A(n535), .B(n445), .ZN(n424) );
  XNOR2_X1 U433 ( .A(G137), .B(G134), .ZN(n445) );
  NAND2_X1 U434 ( .A1(n477), .A2(G214), .ZN(n703) );
  XNOR2_X1 U435 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n473) );
  NAND2_X1 U436 ( .A1(n427), .A2(n660), .ZN(n426) );
  INV_X1 U437 ( .A(G146), .ZN(n490) );
  INV_X1 U438 ( .A(KEYINPUT33), .ZN(n451) );
  INV_X1 U439 ( .A(n672), .ZN(n408) );
  NOR2_X1 U440 ( .A1(n663), .A2(n780), .ZN(n643) );
  XOR2_X1 U441 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n529) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n530) );
  XOR2_X1 U443 ( .A(G122), .B(G107), .Z(n542) );
  XNOR2_X1 U444 ( .A(G134), .B(G116), .ZN(n541) );
  XOR2_X1 U445 ( .A(KEYINPUT106), .B(KEYINPUT9), .Z(n544) );
  INV_X1 U446 ( .A(G237), .ZN(n474) );
  XNOR2_X1 U447 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n522) );
  XNOR2_X1 U448 ( .A(n374), .B(n536), .ZN(n537) );
  INV_X1 U449 ( .A(n615), .ZN(n439) );
  NOR2_X1 U450 ( .A1(n720), .A2(KEYINPUT34), .ZN(n440) );
  INV_X1 U451 ( .A(KEYINPUT92), .ZN(n404) );
  XNOR2_X1 U452 ( .A(n526), .B(n495), .ZN(n738) );
  INV_X1 U453 ( .A(KEYINPUT83), .ZN(n417) );
  INV_X1 U454 ( .A(G902), .ZN(n475) );
  INV_X1 U455 ( .A(n434), .ZN(n727) );
  XNOR2_X1 U456 ( .A(n531), .B(n457), .ZN(n532) );
  XOR2_X1 U457 ( .A(G122), .B(G104), .Z(n534) );
  XNOR2_X1 U458 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n465) );
  XNOR2_X1 U459 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n467) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n480) );
  INV_X1 U461 ( .A(n727), .ZN(n758) );
  XNOR2_X1 U462 ( .A(KEYINPUT16), .B(G122), .ZN(n462) );
  XNOR2_X1 U463 ( .A(G128), .B(G137), .ZN(n498) );
  XNOR2_X1 U464 ( .A(KEYINPUT94), .B(KEYINPUT23), .ZN(n501) );
  XNOR2_X1 U465 ( .A(KEYINPUT108), .B(KEYINPUT105), .ZN(n543) );
  INV_X1 U466 ( .A(KEYINPUT76), .ZN(n433) );
  XOR2_X1 U467 ( .A(G140), .B(KEYINPUT77), .Z(n492) );
  NOR2_X1 U468 ( .A1(n380), .A2(n623), .ZN(n428) );
  XNOR2_X1 U469 ( .A(n450), .B(n612), .ZN(n449) );
  OR2_X1 U470 ( .A1(n611), .A2(n610), .ZN(n450) );
  XNOR2_X1 U471 ( .A(n540), .B(n539), .ZN(n580) );
  INV_X1 U472 ( .A(KEYINPUT86), .ZN(n443) );
  XNOR2_X1 U473 ( .A(n526), .B(n422), .ZN(n657) );
  XNOR2_X1 U474 ( .A(n423), .B(n375), .ZN(n422) );
  NOR2_X1 U475 ( .A1(n421), .A2(n719), .ZN(n642) );
  XNOR2_X1 U476 ( .A(n638), .B(n637), .ZN(n663) );
  NAND2_X1 U477 ( .A1(n636), .A2(n678), .ZN(n638) );
  XNOR2_X1 U478 ( .A(n442), .B(KEYINPUT35), .ZN(n778) );
  NAND2_X1 U479 ( .A1(n438), .A2(n437), .ZN(n442) );
  NAND2_X1 U480 ( .A1(n435), .A2(n440), .ZN(n437) );
  AND2_X1 U481 ( .A1(n580), .A2(n578), .ZN(n674) );
  INV_X1 U482 ( .A(KEYINPUT60), .ZN(n397) );
  XNOR2_X1 U483 ( .A(n740), .B(n739), .ZN(n741) );
  INV_X1 U484 ( .A(KEYINPUT56), .ZN(n395) );
  INV_X1 U485 ( .A(KEYINPUT53), .ZN(n405) );
  AND2_X1 U486 ( .A1(n414), .A2(KEYINPUT2), .ZN(n372) );
  AND2_X1 U487 ( .A1(n477), .A2(G210), .ZN(n373) );
  XOR2_X1 U488 ( .A(n534), .B(n533), .Z(n374) );
  XOR2_X1 U489 ( .A(n522), .B(n521), .Z(n375) );
  AND2_X1 U490 ( .A1(n613), .A2(n632), .ZN(n376) );
  AND2_X1 U491 ( .A1(n723), .A2(n769), .ZN(n378) );
  OR2_X1 U492 ( .A1(n731), .A2(n730), .ZN(n379) );
  NAND2_X1 U493 ( .A1(n365), .A2(n597), .ZN(n380) );
  AND2_X1 U494 ( .A1(n629), .A2(n686), .ZN(n381) );
  AND2_X1 U495 ( .A1(n768), .A2(n728), .ZN(n382) );
  NAND2_X1 U496 ( .A1(n596), .A2(n485), .ZN(n383) );
  AND2_X1 U497 ( .A1(n639), .A2(n691), .ZN(n384) );
  XNOR2_X1 U498 ( .A(n556), .B(KEYINPUT22), .ZN(n385) );
  XOR2_X1 U499 ( .A(n486), .B(KEYINPUT0), .Z(n386) );
  XOR2_X1 U500 ( .A(KEYINPUT66), .B(KEYINPUT19), .Z(n387) );
  XOR2_X1 U501 ( .A(n592), .B(KEYINPUT45), .Z(n388) );
  XNOR2_X1 U502 ( .A(n743), .B(KEYINPUT59), .ZN(n389) );
  XOR2_X1 U503 ( .A(n657), .B(n656), .Z(n390) );
  XOR2_X1 U504 ( .A(n370), .B(n665), .Z(n391) );
  AND2_X1 U505 ( .A1(n728), .A2(KEYINPUT76), .ZN(n392) );
  INV_X1 U506 ( .A(n751), .ZN(n401) );
  NAND2_X1 U507 ( .A1(n429), .A2(n431), .ZN(n393) );
  XNOR2_X1 U508 ( .A(n394), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U509 ( .A1(n400), .A2(n401), .ZN(n394) );
  XNOR2_X1 U510 ( .A(n396), .B(n395), .ZN(G51) );
  NAND2_X1 U511 ( .A1(n399), .A2(n401), .ZN(n396) );
  XNOR2_X1 U512 ( .A(n398), .B(n397), .ZN(G60) );
  NAND2_X1 U513 ( .A1(n402), .A2(n401), .ZN(n398) );
  NAND2_X1 U514 ( .A1(n381), .A2(n448), .ZN(n447) );
  XNOR2_X1 U515 ( .A(n447), .B(n446), .ZN(n427) );
  XNOR2_X1 U516 ( .A(n666), .B(n391), .ZN(n399) );
  XNOR2_X1 U517 ( .A(n658), .B(n390), .ZN(n400) );
  XNOR2_X1 U518 ( .A(n744), .B(n389), .ZN(n402) );
  NAND2_X1 U519 ( .A1(n571), .A2(n384), .ZN(n403) );
  XNOR2_X1 U520 ( .A(n571), .B(n404), .ZN(n577) );
  XNOR2_X2 U521 ( .A(n487), .B(n386), .ZN(n571) );
  XNOR2_X1 U522 ( .A(n444), .B(n443), .ZN(n565) );
  XNOR2_X1 U523 ( .A(n567), .B(n566), .ZN(n781) );
  XNOR2_X1 U524 ( .A(n406), .B(n405), .ZN(G75) );
  NAND2_X1 U525 ( .A1(n416), .A2(n378), .ZN(n406) );
  INV_X1 U526 ( .A(n778), .ZN(n409) );
  XNOR2_X1 U527 ( .A(n410), .B(KEYINPUT87), .ZN(n591) );
  NAND2_X1 U528 ( .A1(n585), .A2(n586), .ZN(n410) );
  NAND2_X1 U529 ( .A1(n419), .A2(n736), .ZN(n418) );
  XNOR2_X1 U530 ( .A(n418), .B(n417), .ZN(n416) );
  INV_X1 U531 ( .A(n758), .ZN(n415) );
  NAND2_X1 U532 ( .A1(n742), .A2(G475), .ZN(n744) );
  INV_X1 U533 ( .A(n655), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n420), .A2(n379), .ZN(n419) );
  INV_X1 U535 ( .A(n732), .ZN(n420) );
  INV_X1 U536 ( .A(n456), .ZN(n421) );
  XNOR2_X1 U537 ( .A(n520), .B(n525), .ZN(n423) );
  NAND2_X2 U538 ( .A1(n425), .A2(n776), .ZN(n768) );
  XNOR2_X2 U539 ( .A(n426), .B(n650), .ZN(n425) );
  NAND2_X1 U540 ( .A1(n369), .A2(n560), .ZN(n444) );
  NAND2_X1 U541 ( .A1(n369), .A2(n428), .ZN(n563) );
  INV_X1 U542 ( .A(n768), .ZN(n429) );
  NAND2_X1 U543 ( .A1(n382), .A2(n432), .ZN(n430) );
  NAND2_X1 U544 ( .A1(n434), .A2(n433), .ZN(n432) );
  XNOR2_X2 U545 ( .A(n593), .B(n388), .ZN(n434) );
  NAND2_X1 U546 ( .A1(n434), .A2(n392), .ZN(n431) );
  INV_X1 U547 ( .A(n577), .ZN(n435) );
  NAND2_X1 U548 ( .A1(n720), .A2(KEYINPUT34), .ZN(n441) );
  XNOR2_X2 U549 ( .A(n488), .B(G131), .ZN(n535) );
  XNOR2_X2 U550 ( .A(G143), .B(G128), .ZN(n550) );
  NAND2_X1 U551 ( .A1(n449), .A2(n376), .ZN(n635) );
  AND2_X1 U552 ( .A1(n449), .A2(n613), .ZN(n633) );
  XNOR2_X2 U553 ( .A(n454), .B(G146), .ZN(n496) );
  NAND2_X1 U554 ( .A1(n455), .A2(n383), .ZN(n487) );
  NAND2_X1 U555 ( .A1(n456), .A2(n455), .ZN(n673) );
  AND2_X1 U556 ( .A1(G214), .A2(n530), .ZN(n457) );
  XOR2_X1 U557 ( .A(KEYINPUT114), .B(n645), .Z(n458) );
  INV_X1 U558 ( .A(KEYINPUT25), .ZN(n511) );
  XNOR2_X1 U559 ( .A(n512), .B(n511), .ZN(n514) );
  XNOR2_X1 U560 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U561 ( .A(n538), .B(n537), .ZN(n743) );
  INV_X1 U562 ( .A(n579), .ZN(n578) );
  XNOR2_X1 U563 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X2 U564 ( .A(KEYINPUT68), .B(G101), .ZN(n524) );
  XNOR2_X1 U565 ( .A(n524), .B(KEYINPUT71), .ZN(n464) );
  XNOR2_X1 U566 ( .A(n752), .B(n464), .ZN(n494) );
  XNOR2_X1 U567 ( .A(n755), .B(n494), .ZN(n472) );
  XNOR2_X1 U568 ( .A(n496), .B(n465), .ZN(n469) );
  NAND2_X1 U569 ( .A1(n769), .A2(G224), .ZN(n466) );
  XNOR2_X1 U570 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U572 ( .A(n470), .B(n489), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n664) );
  XNOR2_X1 U574 ( .A(n473), .B(n475), .ZN(n655) );
  NAND2_X1 U575 ( .A1(n664), .A2(n655), .ZN(n476) );
  NAND2_X1 U576 ( .A1(n475), .A2(n474), .ZN(n477) );
  XNOR2_X2 U577 ( .A(n476), .B(n373), .ZN(n630) );
  NAND2_X1 U578 ( .A1(n630), .A2(n703), .ZN(n479) );
  INV_X1 U579 ( .A(KEYINPUT88), .ZN(n478) );
  XNOR2_X2 U580 ( .A(n479), .B(n478), .ZN(n625) );
  XOR2_X1 U581 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n481) );
  XOR2_X1 U582 ( .A(n481), .B(n480), .Z(n483) );
  NAND2_X1 U583 ( .A1(G952), .A2(n483), .ZN(n718) );
  NOR2_X1 U584 ( .A1(G953), .A2(n718), .ZN(n482) );
  XNOR2_X1 U585 ( .A(n482), .B(KEYINPUT91), .ZN(n596) );
  AND2_X1 U586 ( .A1(n483), .A2(G953), .ZN(n484) );
  NAND2_X1 U587 ( .A1(G902), .A2(n484), .ZN(n594) );
  OR2_X1 U588 ( .A1(n594), .A2(G898), .ZN(n485) );
  INV_X1 U589 ( .A(KEYINPUT67), .ZN(n486) );
  NAND2_X1 U590 ( .A1(G227), .A2(n769), .ZN(n491) );
  XNOR2_X1 U591 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X2 U593 ( .A(n497), .B(KEYINPUT10), .ZN(n767) );
  XOR2_X1 U594 ( .A(G110), .B(G119), .Z(n499) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U596 ( .A(n767), .B(n500), .ZN(n508) );
  XNOR2_X1 U597 ( .A(n501), .B(KEYINPUT93), .ZN(n502) );
  XOR2_X1 U598 ( .A(KEYINPUT24), .B(n502), .Z(n506) );
  NAND2_X1 U599 ( .A1(n769), .A2(G234), .ZN(n504) );
  XNOR2_X1 U600 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n503) );
  XNOR2_X1 U601 ( .A(n504), .B(n503), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G221), .A2(n547), .ZN(n505) );
  XNOR2_X1 U603 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U604 ( .A(n508), .B(n507), .ZN(n748) );
  NOR2_X1 U605 ( .A1(G902), .A2(n748), .ZN(n516) );
  NAND2_X1 U606 ( .A1(n655), .A2(G234), .ZN(n510) );
  XNOR2_X1 U607 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n509) );
  XNOR2_X1 U608 ( .A(n510), .B(n509), .ZN(n517) );
  NAND2_X1 U609 ( .A1(n517), .A2(G217), .ZN(n512) );
  INV_X1 U610 ( .A(KEYINPUT95), .ZN(n513) );
  XNOR2_X2 U611 ( .A(n516), .B(n515), .ZN(n597) );
  AND2_X1 U612 ( .A1(n517), .A2(G221), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n518), .B(KEYINPUT21), .ZN(n691) );
  INV_X1 U614 ( .A(n691), .ZN(n519) );
  NAND2_X1 U615 ( .A1(G210), .A2(n530), .ZN(n521) );
  XNOR2_X1 U616 ( .A(KEYINPUT75), .B(KEYINPUT98), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n693), .B(KEYINPUT6), .ZN(n560) );
  INV_X1 U619 ( .A(n560), .ZN(n623) );
  XNOR2_X1 U620 ( .A(KEYINPUT11), .B(KEYINPUT102), .ZN(n528) );
  XNOR2_X1 U621 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U622 ( .A(n767), .B(n532), .ZN(n538) );
  XNOR2_X1 U623 ( .A(n535), .B(KEYINPUT12), .ZN(n536) );
  NOR2_X1 U624 ( .A1(G902), .A2(n743), .ZN(n540) );
  XOR2_X1 U625 ( .A(KEYINPUT13), .B(G475), .Z(n539) );
  XNOR2_X1 U626 ( .A(n542), .B(n541), .ZN(n546) );
  XNOR2_X1 U627 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U628 ( .A(n546), .B(n545), .Z(n549) );
  NAND2_X1 U629 ( .A1(G217), .A2(n547), .ZN(n548) );
  XNOR2_X1 U630 ( .A(n549), .B(n548), .ZN(n554) );
  XOR2_X1 U631 ( .A(KEYINPUT7), .B(n550), .Z(n552) );
  XOR2_X1 U632 ( .A(KEYINPUT107), .B(KEYINPUT109), .Z(n551) );
  XNOR2_X1 U633 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U634 ( .A(n554), .B(n553), .ZN(n745) );
  NOR2_X1 U635 ( .A1(G902), .A2(n745), .ZN(n555) );
  XNOR2_X1 U636 ( .A(G478), .B(n555), .ZN(n579) );
  OR2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n615) );
  AND2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n639) );
  INV_X1 U639 ( .A(KEYINPUT72), .ZN(n556) );
  INV_X1 U640 ( .A(n597), .ZN(n690) );
  NOR2_X1 U641 ( .A1(n365), .A2(n690), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT113), .ZN(n611) );
  AND2_X1 U643 ( .A1(n558), .A2(n611), .ZN(n559) );
  AND2_X1 U644 ( .A1(n369), .A2(n559), .ZN(n672) );
  XNOR2_X1 U645 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n561), .B(KEYINPUT65), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n587), .A2(KEYINPUT44), .ZN(n586) );
  NOR2_X1 U648 ( .A1(n365), .A2(n597), .ZN(n564) );
  NAND2_X1 U649 ( .A1(n565), .A2(n564), .ZN(n567) );
  INV_X1 U650 ( .A(KEYINPUT112), .ZN(n566) );
  NAND2_X1 U651 ( .A1(n568), .A2(n693), .ZN(n570) );
  INV_X1 U652 ( .A(KEYINPUT100), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n570), .B(n569), .ZN(n698) );
  NAND2_X1 U654 ( .A1(n571), .A2(n698), .ZN(n573) );
  XNOR2_X1 U655 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n572) );
  XNOR2_X1 U656 ( .A(n573), .B(n572), .ZN(n682) );
  NAND2_X1 U657 ( .A1(n688), .A2(n603), .ZN(n574) );
  XNOR2_X1 U658 ( .A(n574), .B(KEYINPUT97), .ZN(n613) );
  INV_X1 U659 ( .A(n693), .ZN(n575) );
  NAND2_X1 U660 ( .A1(n613), .A2(n575), .ZN(n576) );
  OR2_X1 U661 ( .A1(n577), .A2(n576), .ZN(n668) );
  NAND2_X1 U662 ( .A1(n682), .A2(n668), .ZN(n583) );
  XNOR2_X1 U663 ( .A(KEYINPUT110), .B(n674), .ZN(n651) );
  OR2_X1 U664 ( .A1(n580), .A2(n578), .ZN(n680) );
  NOR2_X1 U665 ( .A1(n651), .A2(n678), .ZN(n582) );
  INV_X1 U666 ( .A(KEYINPUT111), .ZN(n581) );
  XNOR2_X1 U667 ( .A(n582), .B(n581), .ZN(n707) );
  INV_X1 U668 ( .A(n707), .ZN(n607) );
  AND2_X1 U669 ( .A1(n583), .A2(n607), .ZN(n584) );
  NOR2_X1 U670 ( .A1(n781), .A2(n584), .ZN(n585) );
  INV_X1 U671 ( .A(n587), .ZN(n589) );
  INV_X1 U672 ( .A(KEYINPUT44), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n593) );
  INV_X1 U675 ( .A(KEYINPUT64), .ZN(n592) );
  INV_X1 U676 ( .A(KEYINPUT2), .ZN(n728) );
  INV_X1 U677 ( .A(n611), .ZN(n600) );
  OR2_X1 U678 ( .A1(n594), .A2(G900), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n631) );
  AND2_X1 U680 ( .A1(n597), .A2(n691), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n631), .A2(n598), .ZN(n622) );
  INV_X1 U682 ( .A(n622), .ZN(n599) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U684 ( .A(KEYINPUT28), .B(KEYINPUT115), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n602), .B(n601), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n607), .A2(n366), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n605), .A2(KEYINPUT80), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n606), .B(KEYINPUT47), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n607), .A2(n673), .ZN(n609) );
  INV_X1 U690 ( .A(KEYINPUT80), .ZN(n608) );
  AND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n618) );
  INV_X1 U692 ( .A(n703), .ZN(n610) );
  INV_X1 U693 ( .A(KEYINPUT30), .ZN(n612) );
  INV_X1 U694 ( .A(n631), .ZN(n614) );
  NOR2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  AND2_X1 U696 ( .A1(n630), .A2(n616), .ZN(n617) );
  AND2_X1 U697 ( .A1(n633), .A2(n617), .ZN(n677) );
  NOR2_X1 U698 ( .A1(n618), .A2(n677), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n621), .B(KEYINPUT73), .ZN(n629) );
  NOR2_X1 U701 ( .A1(n680), .A2(n622), .ZN(n624) );
  AND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n644) );
  NAND2_X1 U703 ( .A1(n644), .A2(n625), .ZN(n627) );
  XNOR2_X1 U704 ( .A(KEYINPUT117), .B(KEYINPUT36), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n628), .A2(n365), .ZN(n686) );
  INV_X1 U707 ( .A(n630), .ZN(n648) );
  XNOR2_X1 U708 ( .A(n648), .B(KEYINPUT38), .ZN(n704) );
  AND2_X1 U709 ( .A1(n704), .A2(n631), .ZN(n632) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(n653) );
  INV_X1 U712 ( .A(n653), .ZN(n636) );
  INV_X1 U713 ( .A(KEYINPUT40), .ZN(n637) );
  INV_X1 U714 ( .A(n639), .ZN(n706) );
  NAND2_X1 U715 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U716 ( .A1(n706), .A2(n708), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT41), .B(n640), .ZN(n719) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n642), .B(n641), .ZN(n780) );
  NAND2_X1 U720 ( .A1(n644), .A2(n703), .ZN(n645) );
  INV_X1 U721 ( .A(n365), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n458), .A2(n646), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n647), .B(KEYINPUT43), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n660) );
  INV_X1 U725 ( .A(KEYINPUT84), .ZN(n650) );
  INV_X1 U726 ( .A(n651), .ZN(n652) );
  OR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT118), .ZN(n776) );
  NAND2_X1 U729 ( .A1(n742), .A2(G472), .ZN(n658) );
  XOR2_X1 U730 ( .A(KEYINPUT119), .B(KEYINPUT62), .Z(n656) );
  INV_X1 U731 ( .A(G952), .ZN(n659) );
  AND2_X1 U732 ( .A1(n659), .A2(G953), .ZN(n751) );
  XNOR2_X1 U733 ( .A(n660), .B(G140), .ZN(G42) );
  XNOR2_X1 U734 ( .A(n661), .B(G119), .ZN(G21) );
  XNOR2_X1 U735 ( .A(G131), .B(KEYINPUT127), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(G33) );
  NAND2_X1 U737 ( .A1(n742), .A2(G210), .ZN(n666) );
  XNOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n665) );
  NOR2_X1 U739 ( .A1(n680), .A2(n668), .ZN(n667) );
  XOR2_X1 U740 ( .A(G104), .B(n667), .Z(G6) );
  INV_X1 U741 ( .A(n674), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n683), .A2(n668), .ZN(n670) );
  XNOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U745 ( .A(G107), .B(n671), .ZN(G9) );
  XOR2_X1 U746 ( .A(G110), .B(n672), .Z(G12) );
  XOR2_X1 U747 ( .A(G128), .B(KEYINPUT29), .Z(n676) );
  NAND2_X1 U748 ( .A1(n366), .A2(n674), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(G30) );
  XOR2_X1 U750 ( .A(G143), .B(n677), .Z(G45) );
  NAND2_X1 U751 ( .A1(n366), .A2(n678), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n679), .B(G146), .ZN(G48) );
  NOR2_X1 U753 ( .A1(n680), .A2(n682), .ZN(n681) );
  XOR2_X1 U754 ( .A(G113), .B(n681), .Z(G15) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U756 ( .A(G116), .B(n684), .Z(G18) );
  XOR2_X1 U757 ( .A(G125), .B(KEYINPUT37), .Z(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(G27) );
  XOR2_X1 U759 ( .A(KEYINPUT51), .B(KEYINPUT122), .Z(n701) );
  NOR2_X1 U760 ( .A1(n688), .A2(n365), .ZN(n689) );
  XNOR2_X1 U761 ( .A(KEYINPUT50), .B(n689), .ZN(n697) );
  NOR2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(n692), .Z(n694) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U765 ( .A(n695), .B(KEYINPUT121), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U769 ( .A1(n719), .A2(n702), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U772 ( .A1(n707), .A2(n708), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n711), .A2(n364), .ZN(n712) );
  XOR2_X1 U775 ( .A(KEYINPUT123), .B(n712), .Z(n713) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U777 ( .A(KEYINPUT52), .B(n715), .Z(n716) );
  XOR2_X1 U778 ( .A(KEYINPUT124), .B(n716), .Z(n717) );
  NOR2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n364), .A2(n719), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n758), .A2(KEYINPUT81), .ZN(n726) );
  NAND2_X1 U783 ( .A1(n768), .A2(KEYINPUT82), .ZN(n724) );
  NAND2_X1 U784 ( .A1(n724), .A2(n728), .ZN(n725) );
  NOR2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n727), .A2(n768), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n728), .A2(KEYINPUT81), .ZN(n729) );
  NAND2_X1 U788 ( .A1(n729), .A2(KEYINPUT82), .ZN(n730) );
  INV_X1 U789 ( .A(KEYINPUT81), .ZN(n733) );
  NOR2_X1 U790 ( .A1(n415), .A2(n733), .ZN(n735) );
  NOR2_X1 U791 ( .A1(n768), .A2(KEYINPUT82), .ZN(n734) );
  NOR2_X1 U792 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U793 ( .A1(n367), .A2(G469), .ZN(n740) );
  XOR2_X1 U794 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n737) );
  NOR2_X1 U795 ( .A1(n751), .A2(n741), .ZN(G54) );
  NAND2_X1 U796 ( .A1(n367), .A2(G478), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n751), .A2(n747), .ZN(G63) );
  NAND2_X1 U799 ( .A1(n367), .A2(G217), .ZN(n749) );
  XNOR2_X1 U800 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U801 ( .A1(n751), .A2(n750), .ZN(G66) );
  XNOR2_X1 U802 ( .A(G101), .B(n752), .ZN(n753) );
  XOR2_X1 U803 ( .A(KEYINPUT126), .B(n753), .Z(n754) );
  XNOR2_X1 U804 ( .A(n368), .B(n754), .ZN(n757) );
  NOR2_X1 U805 ( .A1(G898), .A2(n769), .ZN(n756) );
  NOR2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n765) );
  NAND2_X1 U807 ( .A1(n758), .A2(n769), .ZN(n763) );
  XOR2_X1 U808 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n760) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n759) );
  XNOR2_X1 U810 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U811 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U813 ( .A(n765), .B(n764), .ZN(G69) );
  XOR2_X1 U814 ( .A(n766), .B(n767), .Z(n771) );
  XNOR2_X1 U815 ( .A(n768), .B(n771), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U817 ( .A(n771), .B(G227), .ZN(n772) );
  NAND2_X1 U818 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U819 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U820 ( .A1(n775), .A2(n774), .ZN(G72) );
  XNOR2_X1 U821 ( .A(G134), .B(n776), .ZN(n777) );
  XNOR2_X1 U822 ( .A(n777), .B(KEYINPUT120), .ZN(G36) );
  BUF_X1 U823 ( .A(n778), .Z(n779) );
  XOR2_X1 U824 ( .A(n779), .B(G122), .Z(G24) );
  XOR2_X1 U825 ( .A(G137), .B(n780), .Z(G39) );
  XOR2_X1 U826 ( .A(n371), .B(G101), .Z(G3) );
endmodule

