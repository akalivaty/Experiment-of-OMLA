//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n207), .B2(KEYINPUT2), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(new_n202), .A3(KEYINPUT80), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT80), .B1(new_n211), .B2(new_n202), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216));
  XNOR2_X1  g015(.A(G197gat), .B(G204gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218));
  INV_X1    g017(.A(G211gat), .ZN(new_n219));
  INV_X1    g018(.A(G218gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G211gat), .B(G218gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n217), .A3(new_n221), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n216), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  INV_X1    g029(.A(new_n226), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n223), .B1(new_n221), .B2(new_n217), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n215), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n216), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n230), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT75), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n231), .B2(new_n232), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n225), .A2(KEYINPUT75), .A3(new_n226), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G228gat), .ZN(new_n243));
  INV_X1    g042(.A(G233gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n235), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT86), .ZN(new_n247));
  INV_X1    g046(.A(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT85), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n228), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n216), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n248), .B1(new_n251), .B2(new_n215), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT86), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n242), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n236), .A2(new_n230), .B1(new_n239), .B2(new_n240), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n211), .A2(new_n202), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n258), .A2(new_n212), .B1(new_n204), .B2(new_n209), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n216), .B2(new_n233), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n248), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT84), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(new_n248), .C1(new_n255), .C2(new_n260), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n247), .A2(new_n254), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G50gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G78gat), .ZN(new_n270));
  INV_X1    g069(.A(G106gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n247), .A2(new_n254), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n262), .A2(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n266), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n280), .A2(G22gat), .B1(KEYINPUT88), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT87), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(KEYINPUT88), .A3(G22gat), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n272), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n274), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT70), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G120gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n290), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n290), .B2(new_n298), .ZN(new_n301));
  INV_X1    g100(.A(G134gat), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(new_n295), .B2(new_n297), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT71), .B(KEYINPUT1), .C1(new_n292), .C2(new_n294), .ZN(new_n306));
  OAI21_X1  g105(.A(G127gat), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n298), .A3(new_n299), .ZN(new_n308));
  AOI21_X1  g107(.A(G134gat), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n259), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT4), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n302), .B1(new_n300), .B2(new_n301), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(G134gat), .A3(new_n308), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n315), .A3(new_n259), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n303), .B2(new_n309), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT81), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n320), .A2(new_n236), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n215), .A3(new_n322), .ZN(new_n325));
  AOI211_X1 g124(.A(KEYINPUT82), .B(new_n318), .C1(new_n325), .C2(new_n310), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT5), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n318), .B1(new_n325), .B2(new_n310), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT5), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G85gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  AND4_X1   g135(.A1(KEYINPUT6), .A2(new_n327), .A3(new_n332), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n332), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT6), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n328), .A2(new_n329), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n331), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n342), .A2(KEYINPUT5), .B1(new_n330), .B2(new_n331), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n336), .B(KEYINPUT90), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n337), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT23), .ZN(new_n349));
  NAND2_X1  g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n349), .A2(KEYINPUT68), .A3(new_n352), .A4(new_n350), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT65), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n364), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT66), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n361), .A2(new_n363), .A3(KEYINPUT66), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n361), .A2(new_n362), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT25), .B1(new_n372), .B2(new_n353), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n375));
  AOI21_X1  g174(.A(G190gat), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(KEYINPUT69), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT26), .ZN(new_n382));
  INV_X1    g181(.A(G169gat), .ZN(new_n383));
  INV_X1    g182(.A(G176gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n360), .C1(new_n376), .C2(new_n378), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n373), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n371), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n347), .B1(new_n391), .B2(KEYINPUT29), .ZN(new_n392));
  INV_X1    g191(.A(new_n241), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n360), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n374), .A2(new_n375), .ZN(new_n397));
  INV_X1    g196(.A(G190gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n378), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n361), .A2(new_n362), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(new_n350), .A3(new_n349), .A4(new_n352), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n400), .A2(new_n380), .B1(KEYINPUT25), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n403), .B(new_n404), .C1(new_n358), .C2(new_n370), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT76), .B1(new_n371), .B2(new_n390), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n347), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n395), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI211_X1 g208(.A(KEYINPUT78), .B(new_n347), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n394), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n403), .B1(new_n358), .B2(new_n370), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n408), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT77), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n408), .B1(new_n407), .B2(new_n230), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n241), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT79), .B(new_n394), .C1(new_n409), .C2(new_n410), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT37), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n416), .A2(new_n241), .A3(new_n417), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n409), .A2(new_n410), .ZN(new_n424));
  INV_X1    g223(.A(new_n392), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n241), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n426), .A3(KEYINPUT37), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  XOR2_X1   g227(.A(G8gat), .B(G36gat), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G64gat), .ZN(new_n430));
  INV_X1    g229(.A(G92gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT38), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n413), .A2(new_n418), .A3(new_n419), .A4(new_n433), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n346), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n420), .B(new_n421), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n439), .B2(new_n432), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n288), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n318), .B1(new_n317), .B2(new_n323), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n325), .A2(new_n310), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n318), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT39), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT91), .B(KEYINPUT39), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n344), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n447), .A2(KEYINPUT92), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT92), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(KEYINPUT40), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI221_X1 g253(.A(new_n445), .B1(new_n452), .B2(KEYINPUT40), .C1(new_n449), .C2(new_n450), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n345), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n420), .A2(new_n432), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(KEYINPUT30), .A3(new_n436), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n413), .A2(new_n419), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n418), .A4(new_n433), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT89), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(KEYINPUT89), .A3(new_n461), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n456), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n441), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n337), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n343), .B2(new_n336), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n338), .A2(new_n339), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n288), .B1(new_n472), .B2(new_n462), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n391), .A2(new_n313), .A3(new_n312), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n414), .A2(new_n314), .ZN(new_n476));
  AND2_X1   g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n477), .B(KEYINPUT64), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT72), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT72), .A4(new_n479), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n474), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G71gat), .ZN(new_n488));
  INV_X1    g287(.A(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n484), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n475), .A2(new_n476), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(new_n477), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(KEYINPUT34), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n494), .A2(KEYINPUT34), .B1(new_n495), .B2(new_n478), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI221_X4 g296(.A(new_n474), .B1(new_n485), .B2(new_n490), .C1(new_n482), .C2(new_n483), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n492), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n484), .ZN(new_n500));
  INV_X1    g299(.A(new_n486), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(new_n490), .ZN(new_n502));
  INV_X1    g301(.A(new_n498), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n497), .B1(new_n492), .B2(new_n498), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(new_n503), .A3(new_n496), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT74), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n502), .A2(KEYINPUT74), .A3(new_n503), .A4(new_n496), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT36), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n473), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n512), .ZN(new_n516));
  INV_X1    g315(.A(new_n346), .ZN(new_n517));
  AND4_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n288), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n464), .A2(new_n465), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n288), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n472), .A2(new_n462), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT35), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n467), .A2(new_n514), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT104), .ZN(new_n525));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G71gat), .B(G78gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n529), .B(new_n530), .Z(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(G85gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n532), .B1(new_n533), .B2(new_n431), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT7), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n533), .B2(new_n431), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G99gat), .B(G106gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(KEYINPUT99), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n538), .A2(new_n540), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n540), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n531), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT10), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n529), .B(new_n530), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(new_n544), .A3(new_n542), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n545), .A2(new_n541), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(KEYINPUT102), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT102), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n526), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n384), .ZN(new_n557));
  INV_X1    g356(.A(G204gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n546), .A2(new_n549), .ZN(new_n561));
  INV_X1    g360(.A(new_n526), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n555), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT103), .ZN(new_n565));
  INV_X1    g364(.A(new_n563), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n550), .B2(new_n552), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n525), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n525), .A3(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n524), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G15gat), .B(G22gat), .ZN(new_n574));
  AOI21_X1  g373(.A(G1gat), .B1(new_n574), .B2(KEYINPUT96), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(KEYINPUT96), .A3(G1gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT16), .ZN(new_n578));
  AOI211_X1 g377(.A(new_n575), .B(new_n577), .C1(new_n578), .C2(new_n574), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G8gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT21), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n531), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G183gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n531), .A2(new_n581), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G211gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n590), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n587), .B(new_n593), .Z(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT15), .ZN(new_n598));
  INV_X1    g397(.A(G50gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(G43gat), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(G43gat), .B2(new_n599), .ZN(new_n601));
  INV_X1    g400(.A(G43gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n602), .B2(G50gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n604), .B1(new_n599), .B2(G43gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT94), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n599), .A3(G43gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(KEYINPUT95), .A3(G50gat), .ZN(new_n608));
  AND4_X1   g407(.A1(new_n603), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n601), .B1(new_n609), .B2(KEYINPUT15), .ZN(new_n610));
  INV_X1    g409(.A(G29gat), .ZN(new_n611));
  INV_X1    g410(.A(G36gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT14), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT14), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(G29gat), .B2(G36gat), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n613), .B(new_n615), .C1(new_n611), .C2(new_n612), .ZN(new_n616));
  MUX2_X1   g415(.A(new_n610), .B(new_n601), .S(new_n616), .Z(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n551), .C1(KEYINPUT100), .C2(KEYINPUT17), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(KEYINPUT17), .Z(new_n619));
  AND2_X1   g418(.A1(new_n619), .A2(KEYINPUT100), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n620), .B2(new_n551), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  NAND3_X1  g421(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n597), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n597), .A2(KEYINPUT101), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(KEYINPUT101), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n594), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n619), .A2(new_n580), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n580), .A2(new_n617), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n580), .B(new_n617), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n636), .B(KEYINPUT13), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT11), .B(G169gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G197gat), .ZN(new_n646));
  XOR2_X1   g445(.A(G113gat), .B(G141gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n644), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n573), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n472), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT105), .B(G1gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n519), .ZN(new_n656));
  NAND2_X1  g455(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n578), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n662), .B(new_n663), .C1(new_n658), .C2(new_n656), .ZN(G1325gat));
  INV_X1    g463(.A(new_n652), .ZN(new_n665));
  AOI21_X1  g464(.A(G15gat), .B1(new_n665), .B2(new_n516), .ZN(new_n666));
  INV_X1    g465(.A(new_n507), .ZN(new_n667));
  INV_X1    g466(.A(new_n513), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n666), .B1(G15gat), .B2(new_n671), .ZN(G1326gat));
  NOR2_X1   g471(.A1(new_n652), .A2(new_n288), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NOR2_X1   g474(.A1(new_n524), .A2(new_n632), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n594), .A2(new_n572), .A3(new_n650), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n472), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT45), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n441), .A2(new_n466), .ZN(new_n682));
  INV_X1    g481(.A(new_n288), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n522), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n667), .A3(new_n668), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n520), .A2(new_n523), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n514), .B(KEYINPUT106), .C1(new_n466), .C2(new_n441), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n632), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n524), .B2(new_n632), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(new_n677), .ZN(new_n695));
  INV_X1    g494(.A(new_n472), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n680), .B1(new_n611), .B2(new_n697), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n678), .A2(G36gat), .A3(new_n519), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  INV_X1    g499(.A(new_n519), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT107), .Z(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n703), .B2(new_n612), .ZN(G1329gat));
  INV_X1    g503(.A(new_n516), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n678), .A2(G43gat), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n695), .A2(new_n669), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n708), .A2(KEYINPUT108), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n708), .B2(KEYINPUT108), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT47), .B(new_n707), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n602), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n706), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(KEYINPUT47), .B2(new_n713), .ZN(G1330gat));
  NAND3_X1  g513(.A1(new_n695), .A2(G50gat), .A3(new_n683), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n599), .B1(new_n678), .B2(new_n288), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT48), .ZN(G1331gat));
  XOR2_X1   g517(.A(new_n644), .B(new_n649), .Z(new_n719));
  NOR2_X1   g518(.A1(new_n633), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n689), .A2(new_n572), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n689), .A2(KEYINPUT109), .A3(new_n572), .A4(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n472), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g526(.A1(new_n725), .A2(KEYINPUT110), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n723), .B2(new_n724), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n701), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n734), .ZN(G1333gat));
  NOR3_X1   g534(.A1(new_n725), .A2(G71gat), .A3(new_n705), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n669), .B1(new_n728), .B2(new_n730), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G71gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT50), .ZN(G1334gat));
  OAI21_X1  g538(.A(new_n683), .B1(new_n728), .B2(new_n730), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742));
  INV_X1    g541(.A(new_n594), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n650), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n572), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n694), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g547(.A(KEYINPUT111), .B(new_n746), .C1(new_n692), .C2(new_n693), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n533), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n689), .A2(new_n691), .A3(new_n745), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT51), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n689), .A2(new_n754), .A3(new_n691), .A4(new_n745), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n572), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(new_n472), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n751), .A2(new_n696), .B1(new_n533), .B2(new_n757), .ZN(G1336gat));
  NAND2_X1  g557(.A1(new_n694), .A2(new_n747), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n759), .B2(new_n519), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n519), .A2(G92gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n753), .A2(new_n572), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n746), .B1(new_n692), .B2(new_n693), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n742), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n519), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n769), .B2(new_n431), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n765), .B1(new_n770), .B2(KEYINPUT52), .ZN(new_n771));
  INV_X1    g570(.A(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n701), .B1(new_n748), .B2(new_n749), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(G92gat), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n761), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n764), .B1(new_n771), .B2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n750), .B2(new_n670), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n516), .A2(new_n489), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n756), .B2(new_n778), .ZN(G1338gat));
  NOR3_X1   g578(.A1(new_n756), .A2(G106gat), .A3(new_n288), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n271), .B1(new_n767), .B2(new_n683), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n780), .A2(KEYINPUT53), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n683), .B1(new_n748), .B2(new_n749), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n783), .B2(G106gat), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n550), .A2(new_n562), .A3(new_n552), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n555), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n560), .B1(new_n567), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT55), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n565), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n565), .A2(new_n794), .A3(new_n798), .A4(new_n795), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n639), .A2(new_n649), .A3(new_n642), .A4(new_n643), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n640), .A2(new_n641), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n636), .B1(new_n634), .B2(new_n635), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n648), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n691), .A2(new_n797), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n719), .A2(new_n797), .A3(new_n799), .ZN(new_n806));
  INV_X1    g605(.A(new_n571), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n807), .B2(new_n569), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n787), .B(new_n805), .C1(new_n809), .C2(new_n691), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n691), .B1(new_n806), .B2(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(new_n805), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n743), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n572), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n720), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT115), .B1(new_n817), .B2(new_n288), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n819), .B(new_n683), .C1(new_n814), .C2(new_n816), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n701), .A2(new_n472), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n516), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n650), .ZN(new_n824));
  INV_X1    g623(.A(new_n822), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n521), .B(new_n825), .C1(new_n814), .C2(new_n816), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n293), .A3(new_n719), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(G1340gat));
  NAND4_X1  g627(.A1(new_n821), .A2(new_n572), .A3(new_n516), .A4(new_n822), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n829), .A2(new_n830), .A3(G120gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n829), .B2(G120gat), .ZN(new_n832));
  INV_X1    g631(.A(new_n826), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n572), .A2(new_n291), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT117), .Z(new_n835));
  OAI22_X1  g634(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n835), .ZN(G1341gat));
  AOI21_X1  g635(.A(G127gat), .B1(new_n826), .B2(new_n594), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n823), .A2(new_n299), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n594), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n826), .A2(new_n302), .A3(new_n691), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n823), .B2(new_n632), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(G1343gat));
  OR2_X1    g647(.A1(new_n650), .A2(new_n796), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n691), .B1(new_n849), .B2(new_n808), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n743), .B1(new_n850), .B2(new_n812), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n816), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(KEYINPUT57), .A3(new_n683), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n288), .B1(new_n814), .B2(new_n816), .ZN(new_n854));
  XOR2_X1   g653(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n825), .A2(new_n669), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n650), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n854), .A2(new_n857), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n860), .A2(G141gat), .A3(new_n650), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g662(.A(new_n860), .ZN(new_n864));
  INV_X1    g663(.A(G148gat), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n572), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n854), .A2(new_n855), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n691), .A2(new_n804), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n796), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n850), .A2(new_n870), .A3(KEYINPUT121), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT121), .B1(new_n850), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n743), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n816), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n874), .B2(new_n683), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n815), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n857), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n867), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n867), .B1(new_n858), .B2(new_n815), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n865), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n866), .B1(new_n879), .B2(new_n881), .ZN(G1345gat));
  OAI21_X1  g681(.A(new_n205), .B1(new_n860), .B2(new_n743), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n594), .A2(G155gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n858), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT122), .ZN(G1346gat));
  NOR2_X1   g685(.A1(new_n854), .A2(new_n855), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n888), .B(new_n288), .C1(new_n816), .C2(new_n851), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n691), .B(new_n857), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n856), .A2(KEYINPUT123), .A3(new_n691), .A4(new_n857), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(G162gat), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n864), .A2(new_n206), .A3(new_n691), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(KEYINPUT124), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n519), .A2(new_n696), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n516), .B(new_n901), .C1(new_n818), .C2(new_n820), .ZN(new_n902));
  OAI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n650), .ZN(new_n903));
  AND4_X1   g702(.A1(new_n288), .A2(new_n817), .A3(new_n505), .A4(new_n901), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n383), .A3(new_n719), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n904), .B2(new_n572), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n902), .A2(new_n815), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(G176gat), .ZN(G1349gat));
  NOR2_X1   g708(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n910));
  AND2_X1   g709(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n911));
  OAI21_X1  g710(.A(G183gat), .B1(new_n902), .B2(new_n743), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n904), .A2(new_n397), .A3(new_n594), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AND4_X1   g713(.A1(KEYINPUT125), .A2(new_n912), .A3(KEYINPUT60), .A4(new_n913), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n904), .A2(new_n398), .A3(new_n691), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n902), .A2(new_n632), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(G190gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n918), .B2(G190gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n670), .A2(new_n901), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n876), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(new_n719), .ZN(new_n926));
  INV_X1    g725(.A(new_n924), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n854), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n923), .A3(new_n719), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT126), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n926), .A2(new_n930), .ZN(G1352gat));
  AOI21_X1  g730(.A(new_n558), .B1(new_n877), .B2(new_n927), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n558), .A3(new_n572), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n932), .A2(new_n934), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n219), .A3(new_n594), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n925), .A2(new_n594), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n937), .B2(G211gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n939));
  AOI211_X1 g738(.A(new_n939), .B(new_n219), .C1(new_n925), .C2(new_n594), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n938), .B2(new_n940), .ZN(G1354gat));
  NAND3_X1  g740(.A1(new_n928), .A2(new_n220), .A3(new_n691), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n876), .B2(new_n924), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT127), .B(new_n927), .C1(new_n868), .C2(new_n875), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n944), .A2(new_n691), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n946), .B2(new_n220), .ZN(G1355gat));
endmodule


