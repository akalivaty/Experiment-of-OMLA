//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n193), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n192), .B2(new_n196), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT66), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G143), .B(G146), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n193), .B1(new_n201), .B2(KEYINPUT65), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n216), .A2(new_n208), .A3(new_n210), .A4(new_n211), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n200), .A2(new_n205), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n200), .A2(new_n221), .A3(new_n205), .A4(new_n218), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n208), .A2(new_n210), .A3(new_n213), .A4(new_n211), .ZN(new_n223));
  INV_X1    g037(.A(new_n211), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n207), .A2(G137), .ZN(new_n225));
  OAI21_X1  g039(.A(G131), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n227), .A2(new_n189), .A3(new_n191), .A4(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n190), .B2(G146), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n229), .A2(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n223), .B(new_n226), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n222), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  OR2_X1    g050(.A1(KEYINPUT2), .A2(G113), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n237), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT70), .B1(new_n215), .B2(new_n217), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n202), .A2(new_n203), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n231), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n229), .A2(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n192), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n201), .A2(G128), .A3(new_n229), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n259), .A2(KEYINPUT71), .A3(new_n223), .A4(new_n226), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n253), .A2(KEYINPUT30), .A3(new_n255), .A4(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n234), .A2(new_n247), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n247), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n253), .A2(new_n263), .A3(new_n255), .A4(new_n260), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n266), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT29), .ZN(new_n274));
  INV_X1    g088(.A(new_n231), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n219), .B2(KEYINPUT68), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n263), .B1(new_n276), .B2(new_n222), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n264), .B1(new_n277), .B2(KEYINPUT73), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n232), .A2(KEYINPUT73), .A3(new_n247), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT28), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n253), .A2(new_n231), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n263), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n282), .A2(new_n283), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n280), .A2(new_n272), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n274), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n217), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n290), .A2(new_n248), .A3(new_n250), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n255), .A2(new_n260), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n247), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n264), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT75), .B(new_n247), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n287), .A2(new_n297), .A3(KEYINPUT29), .A4(new_n272), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT76), .B(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n187), .B1(new_n289), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n262), .A2(new_n272), .A3(new_n264), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT31), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n262), .A2(new_n306), .A3(new_n272), .A4(new_n264), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n272), .B1(new_n280), .B2(new_n287), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT32), .B(new_n303), .C1(new_n308), .C2(new_n309), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT77), .A3(new_n313), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n308), .A2(new_n309), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT32), .A4(new_n303), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n302), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT78), .B1(new_n239), .B2(G128), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n319), .A2(KEYINPUT23), .B1(new_n239), .B2(G128), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(KEYINPUT23), .B2(new_n319), .ZN(new_n321));
  XNOR2_X1  g135(.A(G119), .B(G128), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT24), .B(G110), .Z(new_n323));
  OAI22_X1  g137(.A1(new_n321), .A2(G110), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n327), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n329), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n188), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n324), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G140), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n326), .A2(new_n344), .A3(KEYINPUT16), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n332), .B1(new_n345), .B2(KEYINPUT79), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n188), .B1(new_n346), .B2(new_n328), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n333), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n321), .A2(G110), .B1(new_n322), .B2(new_n323), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT80), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT80), .B1(new_n348), .B2(new_n349), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n335), .B(new_n342), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n335), .ZN(new_n354));
  INV_X1    g168(.A(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n341), .B(KEYINPUT83), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n300), .B(new_n353), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n341), .B(KEYINPUT83), .Z(new_n361));
  OAI21_X1  g175(.A(new_n335), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n300), .A4(new_n353), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n300), .B2(G234), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n369), .A3(new_n353), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n318), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G221), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G902), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n290), .A2(new_n248), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT85), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n383), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G104), .B(G107), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n393), .A2(new_n259), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n259), .B1(new_n393), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n378), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n215), .B2(new_n217), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n397), .B2(new_n398), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(KEYINPUT88), .B(new_n402), .C1(new_n397), .C2(new_n398), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n391), .B1(new_n387), .B2(new_n385), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n395), .B1(new_n408), .B2(new_n389), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT10), .B1(new_n409), .B2(new_n259), .ZN(new_n410));
  AND4_X1   g224(.A1(KEYINPUT10), .A2(new_n393), .A3(new_n259), .A4(new_n396), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n387), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n394), .B2(new_n380), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n414), .B2(new_n391), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n389), .B1(new_n388), .B2(new_n392), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(KEYINPUT4), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT87), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n420));
  INV_X1    g234(.A(new_n418), .ZN(new_n421));
  NOR4_X1   g235(.A1(new_n408), .A2(new_n420), .A3(new_n389), .A4(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n251), .B(new_n416), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n378), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n412), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n407), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n337), .A2(G227), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n427), .B(new_n428), .Z(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT84), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n424), .B1(new_n412), .B2(new_n423), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n429), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n426), .A2(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n376), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G469), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n412), .A2(new_n423), .A3(new_n424), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n431), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n407), .A2(new_n425), .A3(new_n429), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(G469), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n300), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n377), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n247), .B(new_n416), .C1(new_n419), .C2(new_n422), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(G113), .C1(KEYINPUT5), .C2(new_n240), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n409), .A2(new_n448), .A3(new_n246), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n446), .A2(new_n451), .A3(new_n449), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n456), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n250), .A2(G125), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(G125), .B2(new_n259), .ZN(new_n459));
  INV_X1    g273(.A(G224), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G953), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n459), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(new_n460), .B2(G953), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n459), .B(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n451), .B(KEYINPUT8), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n448), .A2(new_n246), .ZN(new_n467));
  INV_X1    g281(.A(new_n409), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n469), .B2(new_n449), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n471), .B2(new_n454), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n474), .A3(new_n472), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n445), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n443), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  OR2_X1    g294(.A1(KEYINPUT90), .A2(G143), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT90), .A2(G143), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n481), .A2(new_n482), .B1(new_n267), .B2(G214), .ZN(new_n483));
  INV_X1    g297(.A(G237), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n337), .A3(G214), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT90), .A2(G143), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n482), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n485), .B1(new_n489), .B2(new_n486), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n481), .A2(G214), .A3(new_n267), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n213), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT19), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n330), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n330), .A2(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n188), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n333), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT18), .B(G131), .C1(new_n483), .C2(new_n487), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n330), .B(new_n188), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT18), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n490), .A2(new_n501), .A3(new_n491), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .A4(new_n492), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT91), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n383), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n498), .A2(new_n509), .A3(new_n503), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n488), .A2(new_n492), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT17), .B(G131), .C1(new_n483), .C2(new_n487), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n347), .A3(new_n333), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n507), .A3(new_n503), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n511), .A2(KEYINPUT92), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT92), .B1(new_n511), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n480), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT20), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n480), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n511), .B2(new_n516), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT95), .B1(new_n190), .B2(G128), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n528));
  INV_X1    g342(.A(G128), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(G143), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n190), .A2(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n535), .A3(G134), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n531), .B(new_n532), .C1(new_n534), .C2(new_n207), .ZN(new_n537));
  INV_X1    g351(.A(G122), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G116), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n241), .A2(G122), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n381), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(G107), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT14), .A4(G107), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(KEYINPUT14), .A3(G107), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n531), .A2(new_n207), .A3(new_n532), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n207), .B1(new_n531), .B2(new_n532), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n374), .A2(new_n366), .A3(G953), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n545), .A2(new_n551), .A3(new_n553), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n300), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(G478), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n557), .B(new_n300), .C1(KEYINPUT15), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n515), .A2(new_n503), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n508), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n565), .B2(new_n516), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT94), .B(G475), .Z(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G952), .ZN(new_n570));
  AOI211_X1 g384(.A(G953), .B(new_n570), .C1(G234), .C2(G237), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI211_X1 g386(.A(new_n337), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT21), .B(G898), .Z(new_n575));
  OAI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n526), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n479), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n372), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(new_n389), .ZN(G3));
  OAI21_X1  g394(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n310), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n585));
  INV_X1    g399(.A(new_n371), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n443), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n557), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n556), .A2(KEYINPUT98), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n545), .A2(new_n551), .A3(new_n592), .A4(new_n553), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n552), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n545), .A2(new_n551), .A3(KEYINPUT97), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n554), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT33), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n553), .B1(new_n552), .B2(new_n595), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n588), .B1(new_n601), .B2(new_n597), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n594), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n590), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n561), .B1(new_n605), .B2(new_n300), .ZN(new_n606));
  INV_X1    g420(.A(new_n558), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n561), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT100), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n604), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n603), .B1(new_n602), .B2(new_n594), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n300), .B(new_n589), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G478), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n608), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n568), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n526), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n478), .A2(new_n576), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n443), .A2(new_n586), .ZN(new_n623));
  OAI21_X1  g437(.A(KEYINPUT96), .B1(new_n623), .B2(new_n583), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n587), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n511), .A2(new_n516), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT92), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n511), .A2(new_n516), .A3(KEYINPUT92), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n521), .B1(new_n632), .B2(new_n480), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n521), .B(new_n480), .C1(new_n517), .C2(new_n518), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n618), .A2(new_n563), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n621), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n587), .A2(new_n624), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  OAI21_X1  g455(.A(new_n362), .B1(new_n361), .B2(KEYINPUT36), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n356), .A2(new_n357), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n642), .A2(new_n644), .A3(new_n369), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n365), .B2(new_n367), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n583), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n578), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(new_n637), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n571), .B1(new_n573), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n651), .B(new_n654), .C1(new_n633), .C2(new_n635), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n463), .A2(new_n474), .A3(new_n472), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n474), .B1(new_n463), .B2(new_n472), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n444), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n653), .B(new_n637), .C1(new_n520), .C2(new_n634), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n478), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n659), .A2(new_n662), .A3(new_n443), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n318), .A2(new_n646), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n529), .ZN(G30));
  NAND2_X1  g479(.A1(new_n619), .A2(new_n563), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n646), .A2(new_n444), .ZN(new_n667));
  INV_X1    g481(.A(new_n443), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n653), .B(KEYINPUT39), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n666), .B(new_n667), .C1(new_n670), .C2(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n314), .A2(new_n317), .ZN(new_n672));
  INV_X1    g486(.A(new_n304), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n295), .A2(new_n296), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n271), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n476), .A2(new_n477), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n671), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n302), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n646), .B1(new_n672), .B2(new_n684), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n619), .A2(new_n610), .A3(new_n616), .A4(new_n654), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n479), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  INV_X1    g504(.A(new_n377), .ZN(new_n691));
  INV_X1    g505(.A(G469), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n299), .B1(new_n438), .B2(new_n439), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n442), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT103), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n372), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n622), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n638), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NOR2_X1   g516(.A1(new_n693), .A2(new_n692), .ZN(new_n703));
  INV_X1    g517(.A(new_n441), .ZN(new_n704));
  AOI211_X1 g518(.A(new_n299), .B(new_n704), .C1(new_n438), .C2(new_n439), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n703), .A2(new_n705), .A3(new_n377), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n478), .A2(new_n706), .A3(KEYINPUT104), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n658), .B2(new_n694), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n577), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n685), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NOR2_X1   g526(.A1(new_n621), .A2(new_n666), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n695), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n287), .A2(new_n297), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n271), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n305), .A3(new_n307), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n303), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n582), .A2(new_n586), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND2_X1  g535(.A1(new_n707), .A2(new_n709), .ZN(new_n722));
  AOI221_X4 g536(.A(new_n646), .B1(new_n303), .B2(new_n717), .C1(new_n581), .C2(G472), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n686), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  NAND2_X1  g539(.A1(new_n684), .A2(new_n313), .ZN(new_n726));
  INV_X1    g540(.A(new_n312), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n586), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n476), .A2(new_n444), .A3(new_n477), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n668), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n686), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT42), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n372), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n213), .ZN(G33));
  NAND3_X1  g550(.A1(new_n372), .A2(new_n660), .A3(new_n730), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n692), .B1(new_n433), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n739), .B2(new_n433), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n705), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n691), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n669), .ZN(new_n748));
  INV_X1    g562(.A(new_n729), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n619), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n617), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n755), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT106), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(KEYINPUT106), .A3(new_n758), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n584), .A2(new_n646), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT107), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n750), .B1(new_n765), .B2(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  INV_X1    g581(.A(new_n761), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(new_n759), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n769), .A2(KEYINPUT108), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT108), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n766), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  XNOR2_X1  g588(.A(new_n747), .B(KEYINPUT47), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n318), .A2(new_n371), .A3(new_n686), .A4(new_n749), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NOR2_X1   g594(.A1(new_n729), .A2(new_n694), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n586), .A3(new_n571), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n677), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n620), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(G952), .A3(new_n337), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n572), .B1(new_n757), .B2(new_n758), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n719), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n789), .B2(new_n722), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n781), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n728), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(KEYINPUT48), .B(new_n728), .C1(new_n793), .C2(new_n794), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n790), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT118), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n723), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n680), .A2(new_n444), .A3(new_n694), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT115), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n789), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT50), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n789), .A2(KEYINPUT114), .A3(new_n749), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n703), .A2(new_n705), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n775), .B1(new_n691), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n788), .B2(new_n729), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n807), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n617), .A2(new_n619), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n783), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(KEYINPUT117), .B2(KEYINPUT51), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n805), .B2(KEYINPUT50), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n802), .A2(new_n806), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n818), .A2(new_n822), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n800), .A2(new_n801), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n636), .A2(new_n653), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n685), .A2(new_n569), .A3(new_n826), .A4(new_n730), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n730), .A2(new_n723), .A3(new_n686), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n737), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT111), .ZN(new_n830));
  INV_X1    g644(.A(new_n735), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n625), .A2(new_n648), .A3(new_n720), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n579), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n737), .A2(new_n827), .A3(new_n835), .A4(new_n828), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n478), .A2(new_n526), .A3(new_n576), .A4(new_n651), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT110), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n587), .A2(new_n624), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n837), .A2(KEYINPUT110), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n839), .A2(new_n840), .B1(new_n685), .B2(new_n710), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n372), .B(new_n695), .C1(new_n622), .C2(new_n638), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n834), .A2(new_n836), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n832), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  INV_X1    g659(.A(new_n646), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n479), .A2(new_n666), .A3(new_n846), .A4(new_n653), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n685), .A2(new_n688), .B1(new_n677), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n722), .A2(new_n723), .A3(new_n686), .ZN(new_n849));
  INV_X1    g663(.A(new_n663), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n685), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT112), .B1(new_n664), .B2(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n672), .A2(new_n684), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n846), .A3(new_n850), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n724), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n677), .A2(new_n847), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n858), .A3(new_n689), .A4(new_n859), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n845), .B(new_n853), .C1(KEYINPUT52), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT52), .ZN(new_n862));
  INV_X1    g676(.A(new_n853), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT113), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g678(.A(KEYINPUT53), .B(new_n844), .C1(new_n861), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n834), .A2(new_n841), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n735), .B1(new_n829), .B2(KEYINPUT111), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n836), .A4(new_n842), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n852), .B1(new_n848), .B2(new_n851), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n853), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n866), .A3(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n870), .A2(new_n872), .A3(new_n867), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n844), .B1(new_n861), .B2(new_n864), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n867), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n877), .B2(new_n866), .ZN(new_n878));
  OAI22_X1  g692(.A1(new_n825), .A2(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n371), .A2(new_n445), .A3(new_n377), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n809), .A2(KEYINPUT49), .ZN(new_n883));
  OR4_X1    g697(.A1(new_n680), .A2(new_n752), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n677), .B2(new_n884), .ZN(G75));
  NAND2_X1  g699(.A1(new_n570), .A2(G953), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT120), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n455), .A2(new_n457), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n462), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n873), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n299), .A3(new_n475), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n893), .B(new_n895), .C1(KEYINPUT119), .C2(new_n891), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n888), .B1(new_n897), .B2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n874), .ZN(new_n902));
  INV_X1    g716(.A(new_n892), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n866), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n742), .B(KEYINPUT57), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n440), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n903), .A2(new_n300), .A3(new_n741), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n888), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NOR2_X1   g723(.A1(new_n903), .A2(new_n300), .ZN(new_n910));
  AND2_X1   g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n910), .A2(new_n632), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n632), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n888), .ZN(G60));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n878), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n605), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n902), .A2(new_n904), .A3(new_n605), .A4(new_n917), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n920), .A2(new_n887), .A3(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n892), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n363), .A2(new_n353), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT122), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n892), .A2(new_n644), .A3(new_n642), .A4(new_n925), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n888), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n934), .B(new_n936), .ZN(G66));
  INV_X1    g751(.A(new_n575), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n938), .B2(new_n460), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n868), .A2(new_n842), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n889), .B1(G898), .B2(new_n337), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  AOI21_X1  g758(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n234), .A2(new_n261), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n495), .A2(new_n496), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n670), .A2(new_n729), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n637), .B1(new_n520), .B2(new_n525), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n372), .B(new_n952), .C1(new_n784), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n773), .A2(new_n779), .A3(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n854), .A2(new_n689), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n682), .A3(new_n858), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n951), .B1(new_n959), .B2(G953), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n728), .A2(new_n658), .A3(new_n666), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n748), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n831), .A2(new_n737), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n956), .A2(new_n858), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n773), .A2(new_n779), .A3(new_n337), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n947), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n951), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n957), .B(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n972), .A2(new_n773), .A3(new_n779), .A4(new_n954), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(new_n337), .ZN(new_n974));
  INV_X1    g788(.A(new_n968), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n946), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n960), .A2(new_n947), .A3(new_n968), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT126), .B1(new_n974), .B2(new_n975), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n979), .A3(new_n945), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n273), .B2(new_n673), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n877), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n773), .A2(new_n779), .A3(new_n940), .A4(new_n965), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n265), .A2(new_n271), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n887), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n959), .A2(new_n940), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n983), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n265), .A2(new_n271), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n985), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(G57));
endmodule


