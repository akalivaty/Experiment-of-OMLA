

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G651), .A2(n574), .ZN(n802) );
  XNOR2_X2 U556 ( .A(n595), .B(n594), .ZN(n722) );
  NAND2_X1 U557 ( .A1(n622), .A2(G8), .ZN(n710) );
  XNOR2_X1 U558 ( .A(n597), .B(n596), .ZN(n624) );
  OR2_X1 U559 ( .A1(n685), .A2(n684), .ZN(n689) );
  XNOR2_X1 U560 ( .A(n670), .B(n669), .ZN(n672) );
  NAND2_X1 U561 ( .A1(n668), .A2(n667), .ZN(n670) );
  AND2_X1 U562 ( .A1(n709), .A2(n525), .ZN(n721) );
  INV_X1 U563 ( .A(KEYINPUT93), .ZN(n645) );
  XNOR2_X1 U564 ( .A(n666), .B(n665), .ZN(n683) );
  XNOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT32), .ZN(n690) );
  INV_X1 U566 ( .A(KEYINPUT97), .ZN(n673) );
  NAND2_X1 U567 ( .A1(n754), .A2(n522), .ZN(n756) );
  NOR2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n528) );
  NOR2_X1 U570 ( .A1(n766), .A2(n761), .ZN(n522) );
  XOR2_X1 U571 ( .A(n770), .B(KEYINPUT102), .Z(n523) );
  OR2_X1 U572 ( .A1(n769), .A2(n985), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT89), .B(n708), .ZN(n525) );
  BUF_X1 U574 ( .A(n632), .Z(n652) );
  INV_X1 U575 ( .A(KEYINPUT95), .ZN(n664) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n596) );
  XNOR2_X1 U577 ( .A(n664), .B(KEYINPUT31), .ZN(n665) );
  INV_X1 U578 ( .A(KEYINPUT96), .ZN(n669) );
  INV_X1 U579 ( .A(KEYINPUT84), .ZN(n594) );
  AND2_X1 U580 ( .A1(n695), .A2(n703), .ZN(n696) );
  INV_X1 U581 ( .A(KEYINPUT100), .ZN(n755) );
  INV_X1 U582 ( .A(KEYINPUT17), .ZN(n530) );
  INV_X1 U583 ( .A(G651), .ZN(n553) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n807) );
  NOR2_X2 U585 ( .A1(G2104), .A2(n534), .ZN(n896) );
  NAND2_X1 U586 ( .A1(n899), .A2(G137), .ZN(n532) );
  INV_X1 U587 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U588 ( .A1(n526), .A2(G2104), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT65), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n539), .A2(G101), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(n533) );
  XNOR2_X2 U592 ( .A(n531), .B(n530), .ZN(n899) );
  NAND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n538) );
  INV_X1 U594 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U595 ( .A1(G125), .A2(n896), .ZN(n536) );
  AND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U597 ( .A1(G113), .A2(n895), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X2 U599 ( .A1(n538), .A2(n537), .ZN(G160) );
  NAND2_X1 U600 ( .A1(G138), .A2(n899), .ZN(n541) );
  BUF_X1 U601 ( .A(n539), .Z(n900) );
  NAND2_X1 U602 ( .A1(G102), .A2(n900), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G114), .A2(n895), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G126), .A2(n896), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U607 ( .A1(n545), .A2(n544), .ZN(G164) );
  XOR2_X1 U608 ( .A(G543), .B(KEYINPUT0), .Z(n574) );
  NAND2_X1 U609 ( .A1(n802), .A2(G52), .ZN(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n546), .ZN(n552) );
  NAND2_X1 U611 ( .A1(G90), .A2(n807), .ZN(n548) );
  NOR2_X1 U612 ( .A1(n574), .A2(n553), .ZN(n810) );
  NAND2_X1 U613 ( .A1(G77), .A2(n810), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n557) );
  NOR2_X1 U618 ( .A1(G543), .A2(n553), .ZN(n554) );
  XOR2_X1 U619 ( .A(KEYINPUT1), .B(n554), .Z(n555) );
  XNOR2_X2 U620 ( .A(KEYINPUT66), .B(n555), .ZN(n803) );
  NAND2_X1 U621 ( .A1(G64), .A2(n803), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(G301) );
  INV_X1 U623 ( .A(G301), .ZN(G171) );
  NAND2_X1 U624 ( .A1(n807), .A2(G89), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U626 ( .A1(G76), .A2(n810), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n802), .A2(G51), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G63), .A2(n803), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G88), .A2(n807), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G75), .A2(n810), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n802), .A2(G50), .ZN(n571) );
  NAND2_X1 U639 ( .A1(G62), .A2(n803), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n573), .A2(n572), .ZN(G166) );
  INV_X1 U642 ( .A(G166), .ZN(G303) );
  XOR2_X1 U643 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U644 ( .A1(G87), .A2(n574), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U647 ( .A1(n803), .A2(n577), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n802), .A2(G49), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U650 ( .A1(G73), .A2(n810), .ZN(n580) );
  XNOR2_X1 U651 ( .A(n580), .B(KEYINPUT2), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G48), .A2(n802), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G86), .A2(n807), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n803), .A2(G61), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT82), .B(n583), .Z(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(G305) );
  AND2_X1 U659 ( .A1(G60), .A2(n803), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G47), .A2(n802), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G85), .A2(n807), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n810), .A2(G72), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U666 ( .A1(G40), .A2(G160), .ZN(n595) );
  NOR2_X1 U667 ( .A1(G164), .A2(G1384), .ZN(n724) );
  NAND2_X1 U668 ( .A1(n722), .A2(n724), .ZN(n597) );
  INV_X1 U669 ( .A(n624), .ZN(n621) );
  NAND2_X1 U670 ( .A1(n621), .A2(G1341), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT92), .ZN(n609) );
  NAND2_X1 U672 ( .A1(n803), .A2(G56), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT14), .ZN(n602) );
  NAND2_X1 U674 ( .A1(G43), .A2(n802), .ZN(n600) );
  XOR2_X1 U675 ( .A(KEYINPUT73), .B(n600), .Z(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n807), .A2(G81), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G68), .A2(n810), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT13), .B(n606), .Z(n607) );
  NOR2_X1 U682 ( .A1(n608), .A2(n607), .ZN(n1000) );
  NAND2_X1 U683 ( .A1(n609), .A2(n1000), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n624), .A2(G1996), .ZN(n610) );
  XOR2_X1 U685 ( .A(KEYINPUT26), .B(n610), .Z(n611) );
  NOR2_X2 U686 ( .A1(n612), .A2(n611), .ZN(n629) );
  NAND2_X1 U687 ( .A1(G92), .A2(n807), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n802), .A2(G54), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G66), .A2(n803), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G79), .A2(n810), .ZN(n615) );
  XNOR2_X1 U692 ( .A(KEYINPUT75), .B(n615), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT15), .ZN(n918) );
  NAND2_X1 U696 ( .A1(n629), .A2(n918), .ZN(n628) );
  BUF_X1 U697 ( .A(n621), .Z(n622) );
  NAND2_X1 U698 ( .A1(n622), .A2(G1348), .ZN(n626) );
  INV_X1 U699 ( .A(KEYINPUT91), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n624), .B(n623), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n652), .A2(G2067), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n631) );
  OR2_X1 U704 ( .A1(n918), .A2(n629), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n644) );
  NAND2_X1 U706 ( .A1(n632), .A2(G2072), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT27), .ZN(n635) );
  INV_X1 U708 ( .A(G1956), .ZN(n989) );
  NOR2_X1 U709 ( .A1(n652), .A2(n989), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n647) );
  NAND2_X1 U711 ( .A1(n802), .A2(G53), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n803), .A2(G65), .ZN(n636) );
  XOR2_X1 U713 ( .A(KEYINPUT69), .B(n636), .Z(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G91), .A2(n807), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G78), .A2(n810), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n988) );
  NAND2_X1 U719 ( .A1(n647), .A2(n988), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n650) );
  OR2_X1 U722 ( .A1(n988), .A2(n647), .ZN(n648) );
  XNOR2_X1 U723 ( .A(KEYINPUT28), .B(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT29), .ZN(n656) );
  XOR2_X1 U726 ( .A(G1961), .B(KEYINPUT90), .Z(n950) );
  NAND2_X1 U727 ( .A1(n622), .A2(n950), .ZN(n654) );
  XNOR2_X1 U728 ( .A(KEYINPUT25), .B(G2078), .ZN(n965) );
  NAND2_X1 U729 ( .A1(n652), .A2(n965), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n661) );
  AND2_X1 U731 ( .A1(G171), .A2(n661), .ZN(n655) );
  NOR2_X1 U732 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT94), .ZN(n685) );
  INV_X1 U734 ( .A(n685), .ZN(n668) );
  NOR2_X1 U735 ( .A1(G1966), .A2(n710), .ZN(n671) );
  NOR2_X1 U736 ( .A1(n622), .A2(G2084), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n671), .A2(n675), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT30), .B(n659), .ZN(n660) );
  NOR2_X1 U740 ( .A1(G168), .A2(n660), .ZN(n663) );
  NOR2_X1 U741 ( .A1(G171), .A2(n661), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n666) );
  INV_X1 U743 ( .A(n683), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(n673), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n675), .A2(G8), .ZN(n676) );
  NAND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n713) );
  INV_X1 U748 ( .A(G8), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n622), .A2(G2090), .ZN(n679) );
  NOR2_X1 U750 ( .A1(G1971), .A2(n710), .ZN(n678) );
  NOR2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n680), .A2(G303), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n682), .A2(n681), .ZN(n687) );
  OR2_X1 U754 ( .A1(n683), .A2(n687), .ZN(n684) );
  AND2_X1 U755 ( .A1(G286), .A2(G8), .ZN(n686) );
  OR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(n690), .ZN(n711) );
  NAND2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U760 ( .A(n710), .ZN(n717) );
  NAND2_X1 U761 ( .A1(n987), .A2(n717), .ZN(n699) );
  INV_X1 U762 ( .A(n699), .ZN(n692) );
  AND2_X1 U763 ( .A1(n711), .A2(n692), .ZN(n695) );
  NOR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n698), .A2(KEYINPUT33), .ZN(n693) );
  OR2_X1 U766 ( .A1(n710), .A2(n693), .ZN(n694) );
  XOR2_X1 U767 ( .A(G1981), .B(G305), .Z(n1003) );
  AND2_X1 U768 ( .A1(n694), .A2(n1003), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n713), .A2(n696), .ZN(n705) );
  NOR2_X1 U770 ( .A1(G1971), .A2(G303), .ZN(n697) );
  NOR2_X1 U771 ( .A1(n698), .A2(n697), .ZN(n984) );
  OR2_X1 U772 ( .A1(n699), .A2(n984), .ZN(n701) );
  INV_X1 U773 ( .A(KEYINPUT33), .ZN(n700) );
  NAND2_X1 U774 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U775 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n706) );
  XOR2_X1 U778 ( .A(n706), .B(KEYINPUT24), .Z(n707) );
  NOR2_X1 U779 ( .A1(n710), .A2(n707), .ZN(n708) );
  AND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n719) );
  NOR2_X1 U782 ( .A1(G2090), .A2(G303), .ZN(n714) );
  XOR2_X1 U783 ( .A(KEYINPUT99), .B(n714), .Z(n715) );
  NAND2_X1 U784 ( .A1(G8), .A2(n715), .ZN(n716) );
  OR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n718) );
  AND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n721), .A2(n720), .ZN(n754) );
  INV_X1 U788 ( .A(n722), .ZN(n723) );
  NOR2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U790 ( .A(n725), .B(KEYINPUT85), .Z(n753) );
  INV_X1 U791 ( .A(n753), .ZN(n769) );
  NAND2_X1 U792 ( .A1(G116), .A2(n895), .ZN(n727) );
  NAND2_X1 U793 ( .A1(G128), .A2(n896), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U795 ( .A(n728), .B(KEYINPUT35), .ZN(n734) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(KEYINPUT87), .ZN(n732) );
  NAND2_X1 U797 ( .A1(G140), .A2(n899), .ZN(n730) );
  NAND2_X1 U798 ( .A1(G104), .A2(n900), .ZN(n729) );
  NAND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U800 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U801 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n735), .ZN(n892) );
  XOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .Z(n736) );
  XNOR2_X1 U804 ( .A(KEYINPUT86), .B(n736), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n892), .A2(n758), .ZN(n1027) );
  NOR2_X1 U806 ( .A1(n769), .A2(n1027), .ZN(n766) );
  NAND2_X1 U807 ( .A1(G131), .A2(n899), .ZN(n738) );
  NAND2_X1 U808 ( .A1(G95), .A2(n900), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n742) );
  NAND2_X1 U810 ( .A1(G107), .A2(n895), .ZN(n740) );
  NAND2_X1 U811 ( .A1(G119), .A2(n896), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n741) );
  OR2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n889) );
  NAND2_X1 U814 ( .A1(G1991), .A2(n889), .ZN(n752) );
  NAND2_X1 U815 ( .A1(G141), .A2(n899), .ZN(n749) );
  NAND2_X1 U816 ( .A1(G117), .A2(n895), .ZN(n744) );
  NAND2_X1 U817 ( .A1(G129), .A2(n896), .ZN(n743) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U819 ( .A1(n900), .A2(G105), .ZN(n745) );
  XOR2_X1 U820 ( .A(KEYINPUT38), .B(n745), .Z(n746) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U823 ( .A(n750), .B(KEYINPUT88), .ZN(n890) );
  NAND2_X1 U824 ( .A1(G1996), .A2(n890), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n1030) );
  AND2_X1 U826 ( .A1(n753), .A2(n1030), .ZN(n761) );
  XNOR2_X1 U827 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U828 ( .A(G1986), .B(G290), .Z(n985) );
  NAND2_X1 U829 ( .A1(n757), .A2(n524), .ZN(n771) );
  NOR2_X1 U830 ( .A1(n892), .A2(n758), .ZN(n1019) );
  NOR2_X1 U831 ( .A1(G1996), .A2(n890), .ZN(n1023) );
  NOR2_X1 U832 ( .A1(G1986), .A2(G290), .ZN(n759) );
  NOR2_X1 U833 ( .A1(G1991), .A2(n889), .ZN(n1018) );
  NOR2_X1 U834 ( .A1(n759), .A2(n1018), .ZN(n760) );
  NOR2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U836 ( .A1(n1023), .A2(n762), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n763), .B(KEYINPUT39), .ZN(n764) );
  NOR2_X1 U838 ( .A1(n1019), .A2(n764), .ZN(n765) );
  NOR2_X1 U839 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U840 ( .A(n767), .B(KEYINPUT101), .ZN(n768) );
  NOR2_X1 U841 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U842 ( .A1(n771), .A2(n523), .ZN(n772) );
  XNOR2_X1 U843 ( .A(n772), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U844 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U845 ( .A(G57), .ZN(G237) );
  INV_X1 U846 ( .A(G132), .ZN(G219) );
  INV_X1 U847 ( .A(G82), .ZN(G220) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n773) );
  XNOR2_X1 U849 ( .A(n773), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n775) );
  XNOR2_X1 U851 ( .A(G223), .B(KEYINPUT71), .ZN(n838) );
  NAND2_X1 U852 ( .A1(G567), .A2(n838), .ZN(n774) );
  XNOR2_X1 U853 ( .A(n775), .B(n774), .ZN(G234) );
  NAND2_X1 U854 ( .A1(n1000), .A2(G860), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G301), .A2(G868), .ZN(n776) );
  XNOR2_X1 U856 ( .A(n776), .B(KEYINPUT74), .ZN(n778) );
  INV_X1 U857 ( .A(G868), .ZN(n785) );
  INV_X1 U858 ( .A(n918), .ZN(n992) );
  NAND2_X1 U859 ( .A1(n785), .A2(n992), .ZN(n777) );
  NAND2_X1 U860 ( .A1(n778), .A2(n777), .ZN(G284) );
  XOR2_X1 U861 ( .A(KEYINPUT70), .B(n988), .Z(G299) );
  XNOR2_X1 U862 ( .A(KEYINPUT76), .B(n785), .ZN(n779) );
  NOR2_X1 U863 ( .A1(G286), .A2(n779), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G299), .A2(G868), .ZN(n780) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G297) );
  INV_X1 U866 ( .A(G860), .ZN(n801) );
  NAND2_X1 U867 ( .A1(n801), .A2(G559), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n782), .A2(n918), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT16), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT77), .B(n784), .Z(G148) );
  NAND2_X1 U871 ( .A1(n1000), .A2(n785), .ZN(n786) );
  XOR2_X1 U872 ( .A(KEYINPUT78), .B(n786), .Z(n789) );
  NAND2_X1 U873 ( .A1(G868), .A2(n918), .ZN(n787) );
  NOR2_X1 U874 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U875 ( .A1(n789), .A2(n788), .ZN(G282) );
  NAND2_X1 U876 ( .A1(G123), .A2(n896), .ZN(n790) );
  XOR2_X1 U877 ( .A(KEYINPUT79), .B(n790), .Z(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT18), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G111), .A2(n895), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G135), .A2(n899), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G99), .A2(n900), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n1017) );
  XNOR2_X1 U885 ( .A(n1017), .B(G2096), .ZN(n799) );
  INV_X1 U886 ( .A(G2100), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(G156) );
  NAND2_X1 U888 ( .A1(G559), .A2(n918), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n800), .B(n1000), .ZN(n821) );
  NAND2_X1 U890 ( .A1(n801), .A2(n821), .ZN(n814) );
  NAND2_X1 U891 ( .A1(n802), .A2(G55), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G67), .A2(n803), .ZN(n804) );
  NAND2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT81), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G93), .A2(n807), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n810), .A2(G80), .ZN(n811) );
  XOR2_X1 U898 ( .A(KEYINPUT80), .B(n811), .Z(n812) );
  NOR2_X1 U899 ( .A1(n813), .A2(n812), .ZN(n823) );
  XOR2_X1 U900 ( .A(n814), .B(n823), .Z(G145) );
  XNOR2_X1 U901 ( .A(KEYINPUT83), .B(G305), .ZN(n815) );
  XNOR2_X1 U902 ( .A(n815), .B(G288), .ZN(n816) );
  XNOR2_X1 U903 ( .A(KEYINPUT19), .B(n816), .ZN(n818) );
  XNOR2_X1 U904 ( .A(G290), .B(G166), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n818), .B(n817), .ZN(n820) );
  XOR2_X1 U906 ( .A(n823), .B(G299), .Z(n819) );
  XNOR2_X1 U907 ( .A(n820), .B(n819), .ZN(n921) );
  XNOR2_X1 U908 ( .A(n921), .B(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n822), .A2(G868), .ZN(n825) );
  OR2_X1 U910 ( .A1(G868), .A2(n823), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2084), .A2(G2078), .ZN(n826) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U914 ( .A1(G2090), .A2(n827), .ZN(n828) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U916 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G220), .A2(G219), .ZN(n830) );
  XOR2_X1 U919 ( .A(KEYINPUT22), .B(n830), .Z(n831) );
  NOR2_X1 U920 ( .A1(G218), .A2(n831), .ZN(n832) );
  NAND2_X1 U921 ( .A1(G96), .A2(n832), .ZN(n842) );
  NAND2_X1 U922 ( .A1(n842), .A2(G2106), .ZN(n836) );
  NAND2_X1 U923 ( .A1(G69), .A2(G120), .ZN(n833) );
  NOR2_X1 U924 ( .A1(G237), .A2(n833), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G108), .A2(n834), .ZN(n843) );
  NAND2_X1 U926 ( .A1(n843), .A2(G567), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(n931) );
  NAND2_X1 U928 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U929 ( .A1(n931), .A2(n837), .ZN(n841) );
  NAND2_X1 U930 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(G1996), .B(KEYINPUT106), .ZN(n853) );
  XOR2_X1 U943 ( .A(G1991), .B(G1961), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1966), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G1956), .B(G1971), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1976), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n855) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U956 ( .A(KEYINPUT104), .B(G2067), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2090), .B(G2072), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2096), .B(G2100), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U962 ( .A(G2084), .B(G2078), .Z(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G227) );
  XNOR2_X1 U964 ( .A(G1348), .B(G2454), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(G2430), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(G1341), .ZN(n871) );
  XOR2_X1 U967 ( .A(G2443), .B(G2427), .Z(n867) );
  XNOR2_X1 U968 ( .A(G2438), .B(G2446), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n869) );
  XOR2_X1 U970 ( .A(G2451), .B(G2435), .Z(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n872), .A2(G14), .ZN(n873) );
  XNOR2_X1 U974 ( .A(KEYINPUT103), .B(n873), .ZN(G401) );
  NAND2_X1 U975 ( .A1(G124), .A2(n896), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n895), .A2(G112), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G136), .A2(n899), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G100), .A2(n900), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U982 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G139), .A2(n899), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G103), .A2(n900), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G115), .A2(n895), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G127), .A2(n896), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U990 ( .A1(n887), .A2(n886), .ZN(n1011) );
  XOR2_X1 U991 ( .A(G162), .B(n1011), .Z(n888) );
  XNOR2_X1 U992 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U993 ( .A(n891), .B(n890), .Z(n894) );
  XNOR2_X1 U994 ( .A(G164), .B(n892), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n916) );
  NAND2_X1 U996 ( .A1(G118), .A2(n895), .ZN(n898) );
  NAND2_X1 U997 ( .A1(G130), .A2(n896), .ZN(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT108), .B(KEYINPUT45), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(n899), .A2(G142), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n900), .A2(G106), .ZN(n901) );
  XOR2_X1 U1002 ( .A(KEYINPUT107), .B(n901), .Z(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n914) );
  XOR2_X1 U1006 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n1017), .B(KEYINPUT109), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1009 ( .A(n910), .B(KEYINPUT110), .Z(n912) );
  XNOR2_X1 U1010 ( .A(G160), .B(KEYINPUT111), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n914), .B(n913), .Z(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n917), .ZN(G395) );
  XOR2_X1 U1015 ( .A(n1000), .B(n918), .Z(n920) );
  XNOR2_X1 U1016 ( .A(G286), .B(G171), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n922), .B(n921), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n923), .ZN(G397) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n924), .Z(n927) );
  NOR2_X1 U1022 ( .A1(G401), .A2(n931), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT112), .B(n925), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT113), .B(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(n931), .ZN(G319) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1031 ( .A(G1976), .B(G23), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G22), .B(G1971), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT126), .B(n934), .Z(n936) );
  XNOR2_X1 U1035 ( .A(G1986), .B(G24), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1037 ( .A(KEYINPUT58), .B(n937), .Z(n957) );
  XOR2_X1 U1038 ( .A(G1981), .B(G6), .Z(n938) );
  XNOR2_X1 U1039 ( .A(KEYINPUT121), .B(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(G19), .B(G1341), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT122), .B(n941), .ZN(n946) );
  XOR2_X1 U1043 ( .A(KEYINPUT124), .B(G4), .Z(n943) );
  XNOR2_X1 U1044 ( .A(G1348), .B(KEYINPUT59), .ZN(n942) );
  XNOR2_X1 U1045 ( .A(n943), .B(n942), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(KEYINPUT123), .B(n944), .ZN(n945) );
  NAND2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G20), .B(G1956), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n949), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n950), .B(G5), .ZN(n951) );
  NAND2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(G21), .B(G1966), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1055 ( .A(KEYINPUT125), .B(n955), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n958), .Z(n959) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n959), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(n960), .ZN(n1043) );
  INV_X1 U1060 ( .A(KEYINPUT55), .ZN(n1035) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G35), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1063 ( .A(G26), .B(G2067), .ZN(n961) );
  NOR2_X1 U1064 ( .A1(n962), .A2(n961), .ZN(n970) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n963) );
  NAND2_X1 U1066 ( .A1(n963), .A2(G28), .ZN(n964) );
  XNOR2_X1 U1067 ( .A(n964), .B(KEYINPUT116), .ZN(n968) );
  XOR2_X1 U1068 ( .A(n965), .B(G27), .Z(n966) );
  XNOR2_X1 U1069 ( .A(KEYINPUT118), .B(n966), .ZN(n967) );
  NOR2_X1 U1070 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1072 ( .A(KEYINPUT117), .B(G2072), .Z(n971) );
  XNOR2_X1 U1073 ( .A(G33), .B(n971), .ZN(n972) );
  NOR2_X1 U1074 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1075 ( .A(KEYINPUT53), .B(n974), .ZN(n975) );
  NOR2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1077 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1078 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1079 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1080 ( .A(n1035), .B(n980), .ZN(n982) );
  INV_X1 U1081 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1082 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n983), .ZN(n1041) );
  NAND2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1086 ( .A1(n987), .A2(n986), .ZN(n991) );
  XNOR2_X1 U1087 ( .A(n989), .B(n988), .ZN(n990) );
  NOR2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(G301), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(n992), .B(G1348), .ZN(n993) );
  NOR2_X1 U1091 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1094 ( .A(KEYINPUT120), .B(n999), .Z(n1002) );
  XOR2_X1 U1095 ( .A(n1000), .B(G1341), .Z(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G168), .B(G1966), .ZN(n1004) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(n1005), .B(KEYINPUT57), .ZN(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1101 ( .A(G16), .B(KEYINPUT56), .Z(n1008) );
  XNOR2_X1 U1102 ( .A(KEYINPUT119), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1039) );
  XNOR2_X1 U1104 ( .A(G2072), .B(n1011), .ZN(n1012) );
  XNOR2_X1 U1105 ( .A(n1012), .B(KEYINPUT115), .ZN(n1014) );
  XOR2_X1 U1106 ( .A(G2078), .B(G164), .Z(n1013) );
  NOR2_X1 U1107 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1108 ( .A(KEYINPUT50), .B(n1015), .Z(n1033) );
  XOR2_X1 U1109 ( .A(G160), .B(G2084), .Z(n1016) );
  NOR2_X1 U1110 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(G2090), .B(G162), .Z(n1022) );
  NOR2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1115 ( .A(n1024), .B(KEYINPUT51), .ZN(n1025) );
  NOR2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1119 ( .A(KEYINPUT114), .B(n1031), .Z(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1121 ( .A(KEYINPUT52), .B(n1034), .ZN(n1036) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(G29), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1126 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1127 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1128 ( .A(G311), .ZN(G150) );
endmodule

