//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033, new_n1034, new_n1035;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT13), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G1gat), .B2(new_n204), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G8gat), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n210), .C1(G1gat), .C2(new_n204), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n209), .A2(KEYINPUT93), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT93), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G43gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(KEYINPUT90), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n226), .A2(new_n227), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n216), .B(new_n218), .C1(KEYINPUT90), .C2(KEYINPUT15), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n222), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT91), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  OR3_X1    g031(.A1(new_n228), .A2(new_n221), .A3(new_n219), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n232), .B(new_n233), .C1(new_n212), .C2(new_n213), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n203), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(KEYINPUT17), .A3(new_n233), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n209), .A2(new_n211), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(new_n232), .B2(new_n233), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n235), .B(new_n202), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n240), .A2(new_n242), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n235), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  INV_X1    g047(.A(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT11), .B(G169gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT12), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n245), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n245), .B2(new_n247), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G120gat), .B(G148gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(G176gat), .B(G204gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(KEYINPUT95), .A2(G57gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G64gat), .ZN(new_n261));
  INV_X1    g060(.A(G71gat), .ZN(new_n262));
  INV_X1    g061(.A(G78gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT9), .ZN(new_n264));
  NAND2_X1  g063(.A1(G71gat), .A2(G78gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT96), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT96), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n261), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT94), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT94), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(G71gat), .B2(G78gat), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n271), .A2(new_n273), .A3(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(G64gat), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n275), .A2(G57gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(G57gat), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT9), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n268), .A2(new_n270), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G99gat), .A2(G106gat), .ZN(new_n280));
  INV_X1    g079(.A(G85gat), .ZN(new_n281));
  INV_X1    g080(.A(G92gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(KEYINPUT8), .A2(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n281), .B2(new_n282), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G99gat), .B(G106gat), .Z(new_n288));
  AND2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n279), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n278), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n261), .A2(new_n269), .A3(new_n266), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n269), .B1(new_n261), .B2(new_n266), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n287), .B(new_n288), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(KEYINPUT99), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT99), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT10), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT10), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n292), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G230gat), .ZN(new_n305));
  INV_X1    g104(.A(G233gat), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n302), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n308), .A3(new_n301), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT100), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n309), .A2(new_n310), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n259), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n259), .ZN(new_n317));
  AOI211_X1 g116(.A(new_n317), .B(new_n314), .C1(new_n307), .C2(new_n312), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n256), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT21), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n212), .A2(new_n213), .B1(new_n321), .B2(new_n296), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n322), .B(KEYINPUT98), .Z(new_n323));
  AND2_X1   g122(.A1(G231gat), .A2(G233gat), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n279), .A2(KEYINPUT21), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n325), .B(new_n326), .C1(KEYINPUT21), .C2(new_n279), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n332));
  XNOR2_X1  g131(.A(G183gat), .B(G211gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G155gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT20), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n334), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n329), .A2(new_n337), .A3(new_n330), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n234), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n238), .B(new_n297), .C1(new_n343), .C2(new_n241), .ZN(new_n344));
  XOR2_X1   g143(.A(G134gat), .B(G162gat), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(G232gat), .A2(G233gat), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n234), .A2(new_n291), .B1(KEYINPUT41), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n344), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n346), .B1(new_n344), .B2(new_n348), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n347), .A2(KEYINPUT41), .ZN(new_n351));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR3_X1    g153(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n349), .B2(new_n350), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(new_n281), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT0), .B(G57gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT81), .A2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT2), .ZN(new_n365));
  INV_X1    g164(.A(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G162gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(G141gat), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(KEYINPUT80), .ZN(new_n374));
  OAI21_X1  g173(.A(G148gat), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G148gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G141gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(G148gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT79), .A2(KEYINPUT2), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n378), .A2(KEYINPUT3), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n373), .A2(KEYINPUT80), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n371), .A2(G141gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n376), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n377), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n365), .B(new_n379), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n381), .A2(new_n384), .ZN(new_n393));
  INV_X1    g192(.A(new_n379), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G127gat), .B(G134gat), .ZN(new_n398));
  XOR2_X1   g197(.A(G113gat), .B(G120gat), .Z(new_n399));
  INV_X1    g198(.A(KEYINPUT1), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n400), .ZN(new_n402));
  INV_X1    g201(.A(G120gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT68), .ZN(new_n405));
  INV_X1    g204(.A(G113gat), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(G120gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(G120gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT69), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n402), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT69), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT82), .B(new_n401), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n410), .ZN(new_n415));
  INV_X1    g214(.A(new_n402), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n401), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n397), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n397), .B(KEYINPUT83), .C1(new_n413), .C2(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n392), .A2(new_n395), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n426), .A2(KEYINPUT4), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n401), .B1(new_n411), .B2(new_n412), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n375), .A2(new_n377), .ZN(new_n431));
  INV_X1    g230(.A(new_n370), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n385), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n424), .A2(KEYINPUT5), .A3(new_n425), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n428), .A2(new_n434), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n422), .B2(new_n423), .ZN(new_n439));
  INV_X1    g238(.A(new_n425), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n426), .A2(KEYINPUT82), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n430), .A2(new_n414), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n433), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n426), .A2(new_n427), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n439), .A2(new_n425), .B1(KEYINPUT5), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n363), .B1(new_n437), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n442), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT83), .B1(new_n449), .B2(new_n397), .ZN(new_n450));
  INV_X1    g249(.A(new_n423), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n425), .B(new_n435), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n362), .A3(new_n436), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n437), .A2(new_n446), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT6), .A4(new_n362), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n362), .A4(new_n436), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G64gat), .B(G92gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT77), .ZN(new_n464));
  XNOR2_X1  g263(.A(G8gat), .B(G36gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n466), .B(KEYINPUT78), .Z(new_n467));
  XOR2_X1   g266(.A(G197gat), .B(G204gat), .Z(new_n468));
  NOR2_X1   g267(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(G218gat), .A3(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT73), .B(KEYINPUT22), .Z(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G211gat), .B(G218gat), .Z(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT75), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G197gat), .B(G204gat), .ZN(new_n478));
  AND2_X1   g277(.A1(KEYINPUT74), .A2(G211gat), .ZN(new_n479));
  INV_X1    g278(.A(G218gat), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n479), .A2(new_n469), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n475), .A2(KEYINPUT75), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G226gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(G169gat), .ZN(new_n488));
  INV_X1    g287(.A(G176gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT64), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(G169gat), .B2(G176gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT26), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT67), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT26), .B1(new_n490), .B2(new_n492), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G169gat), .A2(G176gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(G169gat), .A2(G176gat), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(new_n494), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n496), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G190gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n506));
  AND2_X1   g305(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G183gat), .A2(G190gat), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n512));
  AOI21_X1  g311(.A(G190gat), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n509), .B(new_n510), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n520));
  INV_X1    g319(.A(G183gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n501), .A2(KEYINPUT23), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G169gat), .B2(G176gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n527), .A3(new_n500), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n517), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(KEYINPUT65), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT65), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n531), .A3(new_n518), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n530), .A2(new_n520), .A3(new_n522), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n493), .A2(KEYINPUT23), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(KEYINPUT25), .A3(new_n500), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n504), .A2(new_n516), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n487), .B1(new_n538), .B2(KEYINPUT29), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n513), .A2(new_n514), .ZN(new_n540));
  INV_X1    g339(.A(new_n510), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n513), .B2(new_n506), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n503), .B1(new_n497), .B2(new_n498), .ZN(new_n543));
  AOI211_X1 g342(.A(KEYINPUT67), .B(KEYINPUT26), .C1(new_n490), .C2(new_n492), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n540), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n529), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n487), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT76), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n550));
  AOI211_X1 g349(.A(new_n550), .B(new_n487), .C1(new_n545), .C2(new_n546), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n486), .B(new_n539), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n477), .A2(new_n485), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n487), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n467), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(new_n557), .A3(new_n466), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT30), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(KEYINPUT30), .B2(new_n559), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n462), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT85), .ZN(new_n564));
  XNOR2_X1  g363(.A(G211gat), .B(G218gat), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT29), .B1(new_n483), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n474), .A2(new_n475), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT3), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT29), .B1(new_n433), .B2(new_n387), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n568), .A2(new_n433), .B1(new_n569), .B2(new_n486), .ZN(new_n570));
  NAND2_X1  g369(.A1(G228gat), .A2(G233gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n554), .B1(new_n427), .B2(KEYINPUT3), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(new_n553), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT29), .B1(new_n477), .B2(new_n485), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n427), .B1(new_n574), .B2(KEYINPUT3), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G22gat), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n564), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G78gat), .B(G106gat), .Z(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT31), .B(G50gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT86), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n573), .A2(new_n575), .ZN(new_n584));
  INV_X1    g383(.A(new_n571), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n554), .B1(new_n474), .B2(new_n475), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n483), .A2(new_n565), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n387), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n588), .A2(new_n427), .B1(new_n572), .B2(new_n553), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n584), .B(new_n577), .C1(new_n585), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT85), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n581), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n486), .A2(new_n554), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n433), .B1(new_n594), .B2(new_n387), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n585), .B1(new_n569), .B2(new_n486), .ZN(new_n596));
  OAI22_X1  g395(.A1(new_n589), .A2(new_n585), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G22gat), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(new_n590), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n583), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n583), .B2(new_n593), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G227gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n502), .B1(new_n495), .B2(KEYINPUT67), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n515), .B1(new_n605), .B2(new_n499), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n535), .B1(KEYINPUT23), .B2(new_n493), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n523), .A2(new_n525), .A3(new_n527), .A4(new_n500), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n533), .B1(new_n608), .B2(new_n517), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n426), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n430), .A2(new_n545), .A3(new_n546), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n611), .B1(new_n538), .B2(new_n430), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT32), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G15gat), .B(G43gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G99gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND3_X1  g420(.A1(new_n616), .A2(new_n618), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT70), .B1(new_n547), .B2(new_n426), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(new_n603), .A3(new_n610), .A4(new_n612), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT34), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n621), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n615), .B(KEYINPUT32), .C1(new_n617), .C2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT71), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n622), .B2(new_n628), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI211_X1 g431(.A(KEYINPUT71), .B(new_n626), .C1(new_n628), .C2(new_n622), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n602), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT35), .B1(new_n563), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n622), .A2(new_n628), .ZN(new_n636));
  INV_X1    g435(.A(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(KEYINPUT72), .A3(new_n629), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT72), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT35), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n462), .A3(new_n642), .A4(new_n562), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n598), .A2(new_n590), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n592), .B1(new_n591), .B2(new_n581), .ZN(new_n646));
  AOI211_X1 g445(.A(KEYINPUT86), .B(new_n582), .C1(new_n590), .C2(KEYINPUT85), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n583), .A2(new_n593), .A3(new_n599), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n563), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n439), .A2(new_n425), .A3(new_n652), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n443), .A2(new_n440), .A3(new_n444), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT39), .B(new_n654), .C1(new_n439), .C2(new_n425), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n655), .A3(new_n363), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n653), .A2(new_n655), .A3(KEYINPUT40), .A4(new_n363), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n658), .A2(new_n561), .A3(new_n455), .A4(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n466), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n547), .A2(new_n548), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n486), .B1(new_n539), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n550), .B1(new_n538), .B2(new_n487), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n548), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n555), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n666), .B2(new_n486), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT37), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT89), .B(new_n661), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT89), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n552), .B2(new_n557), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n466), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT88), .B(KEYINPUT38), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n666), .A2(new_n553), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n539), .A2(new_n662), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n668), .B1(new_n678), .B2(new_n486), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n675), .B(new_n467), .C1(new_n677), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n559), .B1(new_n680), .B2(new_n673), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n602), .B(new_n660), .C1(new_n462), .C2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT36), .B1(new_n632), .B2(new_n633), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n639), .A2(new_n640), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n651), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n320), .B(new_n358), .C1(new_n644), .C2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n462), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g491(.A1(new_n689), .A2(new_n561), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(KEYINPUT42), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT101), .Z(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n693), .B2(new_n210), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(G1325gat));
  AOI21_X1  g499(.A(G15gat), .B1(new_n689), .B2(new_n641), .ZN(new_n701));
  INV_X1    g500(.A(new_n687), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(G15gat), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n689), .B2(new_n703), .ZN(G1326gat));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n650), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n577), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  AOI21_X1  g507(.A(new_n357), .B1(new_n644), .B2(new_n688), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n635), .A2(KEYINPUT103), .A3(new_n643), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT103), .B1(new_n635), .B2(new_n643), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n688), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n357), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n342), .A2(new_n320), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n462), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n709), .A2(new_n718), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n224), .A3(new_n690), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n225), .A3(new_n561), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n719), .B2(new_n562), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(G1329gat));
  AOI21_X1  g530(.A(G43gat), .B1(new_n639), .B2(new_n640), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n709), .A2(new_n718), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n709), .A2(KEYINPUT105), .A3(new_n718), .A4(new_n732), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n651), .A2(new_n683), .A3(new_n687), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT35), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n460), .B(new_n458), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n561), .B1(new_n741), .B2(new_n456), .ZN(new_n742));
  INV_X1    g541(.A(new_n633), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n638), .A2(KEYINPUT71), .A3(new_n629), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n650), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n740), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  AND4_X1   g545(.A1(new_n462), .A2(new_n641), .A3(new_n642), .A4(new_n562), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n635), .A2(KEYINPUT103), .A3(new_n643), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n738), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n716), .B1(new_n750), .B2(new_n357), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(new_n702), .A3(new_n718), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n737), .B1(new_n753), .B2(G43gat), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(KEYINPUT106), .A3(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(KEYINPUT106), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n754), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n756), .A2(new_n759), .ZN(G1330gat));
  NAND4_X1  g559(.A1(new_n751), .A2(new_n650), .A3(new_n718), .A4(new_n752), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G50gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n602), .A2(G50gat), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n721), .A2(new_n763), .B1(KEYINPUT107), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n764), .A2(KEYINPUT107), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1331gat));
  OR2_X1    g567(.A1(new_n316), .A2(new_n318), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n342), .A2(new_n769), .A3(new_n357), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n750), .A2(new_n256), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n690), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n561), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT49), .B(G64gat), .Z(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1333gat));
  AOI21_X1  g576(.A(new_n262), .B1(new_n771), .B2(new_n702), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n641), .B(KEYINPUT108), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(G71gat), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n778), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n771), .A2(new_n650), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n342), .B2(new_n256), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n254), .A2(new_n255), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n341), .A2(KEYINPUT109), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n713), .A2(new_n714), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n748), .A2(new_n749), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n357), .B1(new_n793), .B2(new_n688), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT51), .A3(new_n789), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n319), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n281), .A3(new_n690), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n319), .B1(new_n786), .B2(new_n788), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n717), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(new_n690), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n797), .B1(new_n800), .B2(new_n281), .ZN(G1336gat));
  NAND4_X1  g600(.A1(new_n717), .A2(KEYINPUT110), .A3(new_n561), .A4(new_n798), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n751), .A2(new_n561), .A3(new_n752), .A4(new_n798), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n805), .A3(G92gat), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n562), .A2(G92gat), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n794), .B2(new_n789), .ZN(new_n810));
  AND4_X1   g609(.A1(KEYINPUT51), .A2(new_n713), .A3(new_n714), .A4(new_n789), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n769), .B(new_n807), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n803), .A2(G92gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n815), .ZN(G1337gat));
  AND2_X1   g615(.A1(new_n799), .A2(new_n702), .ZN(new_n817));
  INV_X1    g616(.A(G99gat), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n810), .A2(new_n811), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n641), .A2(new_n818), .A3(new_n769), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT111), .Z(new_n821));
  OAI22_X1  g620(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(new_n821), .ZN(G1338gat));
  NOR2_X1   g621(.A1(new_n602), .A2(G106gat), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n769), .B(new_n823), .C1(new_n810), .C2(new_n811), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n751), .A2(new_n650), .A3(new_n752), .A4(new_n798), .ZN(new_n825));
  XNOR2_X1  g624(.A(KEYINPUT112), .B(G106gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1339gat));
  NAND2_X1  g631(.A1(new_n743), .A2(new_n744), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  INV_X1    g633(.A(new_n298), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT99), .B1(new_n296), .B2(new_n297), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n301), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n303), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n304), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n308), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n307), .A3(KEYINPUT54), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  OAI221_X1 g642(.A(new_n843), .B1(new_n305), .B2(new_n306), .C1(new_n302), .C2(new_n304), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n259), .A4(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n308), .B1(new_n839), .B2(new_n840), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n315), .B1(new_n846), .B2(new_n311), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n317), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n317), .B1(new_n846), .B2(new_n843), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT55), .B1(new_n850), .B2(new_n842), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n834), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n841), .A2(new_n307), .A3(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n844), .A2(new_n259), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n856), .A2(KEYINPUT113), .A3(new_n848), .A4(new_n845), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n787), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n202), .B1(new_n246), .B2(new_n235), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n235), .A2(new_n236), .A3(new_n203), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n252), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n245), .A2(new_n247), .A3(new_n253), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n769), .A2(new_n864), .A3(KEYINPUT114), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n319), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n357), .B1(new_n858), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(new_n355), .A3(new_n356), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n852), .B2(new_n857), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n342), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NOR4_X1   g672(.A1(new_n341), .A2(new_n256), .A3(new_n769), .A4(new_n714), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n602), .B(new_n833), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n462), .A2(new_n561), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n406), .A3(new_n256), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n641), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n602), .B1(new_n873), .B2(new_n874), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT115), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n883), .B(new_n602), .C1(new_n873), .C2(new_n874), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n406), .B1(new_n885), .B2(new_n256), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n879), .B1(new_n888), .B2(new_n889), .ZN(G1340gat));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(new_n884), .ZN(new_n892));
  INV_X1    g691(.A(new_n880), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(new_n769), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G120gat), .ZN(new_n895));
  NOR4_X1   g694(.A1(new_n875), .A2(G120gat), .A3(new_n319), .A4(new_n877), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT117), .B(new_n896), .C1(new_n894), .C2(G120gat), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1341gat));
  AOI21_X1  g699(.A(G127gat), .B1(new_n878), .B2(new_n342), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n342), .A2(G127gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(new_n885), .B2(new_n902), .ZN(G1342gat));
  NAND2_X1  g702(.A1(new_n714), .A2(new_n562), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n875), .A2(G134gat), .A3(new_n462), .A4(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n714), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G134gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1343gat));
  XNOR2_X1  g708(.A(KEYINPUT80), .B(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n650), .C1(new_n873), .C2(new_n874), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n702), .A2(new_n877), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT118), .B1(new_n854), .B2(new_n855), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n850), .A2(new_n916), .A3(new_n842), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n853), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n845), .A2(new_n848), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n256), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n769), .A2(new_n864), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n714), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n341), .B1(new_n922), .B2(new_n871), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n874), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n341), .C1(new_n922), .C2(new_n871), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n602), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n912), .B(new_n913), .C1(new_n926), .C2(new_n911), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n910), .B1(new_n927), .B2(new_n787), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(KEYINPUT58), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n869), .A2(new_n872), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n341), .ZN(new_n933));
  INV_X1    g732(.A(new_n874), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n650), .A3(new_n913), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n787), .A2(G141gat), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n937), .A2(new_n938), .B1(new_n929), .B2(KEYINPUT58), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n928), .A2(new_n931), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n931), .B1(new_n928), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1344gat));
  NOR3_X1   g741(.A1(new_n936), .A2(G148gat), .A3(new_n319), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n650), .B1(new_n873), .B2(new_n874), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n602), .A2(KEYINPUT57), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n714), .A2(new_n919), .A3(new_n864), .A4(new_n856), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n922), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n787), .A2(new_n849), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n953), .A2(new_n918), .B1(new_n769), .B2(new_n864), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n952), .B(new_n949), .C1(new_n954), .C2(new_n714), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n951), .A2(new_n341), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n948), .B1(new_n956), .B2(new_n874), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n947), .A2(new_n957), .A3(new_n769), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n913), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n945), .B1(new_n959), .B2(G148gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n927), .A2(new_n319), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n945), .A2(G148gat), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n944), .B1(new_n960), .B2(new_n963), .ZN(G1345gat));
  OAI21_X1  g763(.A(new_n368), .B1(new_n936), .B2(new_n341), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n342), .A2(G155gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n927), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n967), .B(new_n968), .ZN(G1346gat));
  XNOR2_X1  g768(.A(KEYINPUT81), .B(G162gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n927), .B2(new_n357), .ZN(new_n971));
  OR4_X1    g770(.A1(new_n970), .A2(new_n702), .A3(new_n462), .A4(new_n904), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n946), .B2(new_n972), .ZN(G1347gat));
  NOR2_X1   g772(.A1(new_n690), .A2(new_n562), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n875), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(new_n488), .A3(new_n256), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n975), .A2(new_n779), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n882), .B2(new_n884), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n979), .A2(new_n256), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n980), .B2(new_n488), .ZN(G1348gat));
  AOI21_X1  g780(.A(G176gat), .B1(new_n976), .B2(new_n769), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n319), .A2(new_n489), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n979), .B2(new_n983), .ZN(G1349gat));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n985), .A2(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n521), .B1(new_n979), .B2(new_n342), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n341), .B1(new_n511), .B2(new_n512), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n976), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n985), .A2(KEYINPUT60), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n986), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n986), .ZN(new_n993));
  AOI22_X1  g792(.A1(new_n976), .A2(new_n988), .B1(new_n985), .B2(KEYINPUT60), .ZN(new_n994));
  AOI211_X1 g793(.A(new_n341), .B(new_n978), .C1(new_n882), .C2(new_n884), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n993), .B(new_n994), .C1(new_n995), .C2(new_n521), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n992), .A2(new_n996), .ZN(G1350gat));
  NAND3_X1  g796(.A1(new_n976), .A2(new_n505), .A3(new_n714), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n979), .A2(new_n714), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(G190gat), .ZN(new_n1001));
  AOI211_X1 g800(.A(KEYINPUT61), .B(new_n505), .C1(new_n979), .C2(new_n714), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(G1351gat));
  AND2_X1   g802(.A1(new_n947), .A2(new_n957), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n975), .A2(new_n702), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1004), .A2(new_n256), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G197gat), .ZN(new_n1007));
  INV_X1    g806(.A(new_n946), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(new_n1005), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1010), .A2(new_n249), .A3(new_n256), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1007), .A2(new_n1011), .ZN(G1352gat));
  OR2_X1    g811(.A1(new_n319), .A2(G204gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(KEYINPUT62), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n1009), .A2(KEYINPUT62), .A3(new_n1013), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n958), .A2(new_n1005), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1017), .B1(new_n1018), .B2(G204gat), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1019), .ZN(G1353gat));
  NAND4_X1  g819(.A1(new_n947), .A2(new_n957), .A3(new_n342), .A4(new_n1005), .ZN(new_n1021));
  NAND3_X1  g820(.A1(new_n1021), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1021), .A2(G211gat), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT63), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g826(.A1(new_n1021), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI211_X1 g828(.A(new_n1010), .B(new_n342), .C1(new_n469), .C2(new_n479), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1029), .A2(new_n1030), .ZN(G1354gat));
  NAND2_X1  g830(.A1(new_n714), .A2(G218gat), .ZN(new_n1032));
  XNOR2_X1  g831(.A(new_n1032), .B(KEYINPUT127), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n1004), .A2(new_n1005), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n480), .B1(new_n1009), .B2(new_n357), .ZN(new_n1035));
  AND2_X1   g834(.A1(new_n1034), .A2(new_n1035), .ZN(G1355gat));
endmodule


