//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G143), .B1(new_n191), .B2(G214), .ZN(new_n194));
  OAI21_X1  g008(.A(G131), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(new_n192), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT16), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT75), .A2(G125), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT75), .A2(G125), .ZN(new_n204));
  OAI21_X1  g018(.A(G140), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(G125), .A2(G140), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n202), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT75), .A2(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT75), .A2(G125), .ZN(new_n210));
  AOI211_X1 g024(.A(KEYINPUT16), .B(G140), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n201), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  INV_X1    g027(.A(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n202), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n213), .B2(G140), .ZN(new_n216));
  OAI211_X1 g030(.A(G146), .B(new_n215), .C1(new_n216), .C2(new_n202), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n196), .A2(new_n192), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT17), .A3(G131), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n200), .A2(new_n212), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G113), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(G146), .ZN(new_n224));
  XNOR2_X1  g038(.A(G125), .B(G140), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n201), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT18), .A2(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n196), .A2(new_n192), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n218), .A2(KEYINPUT18), .A3(G131), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n220), .A2(new_n223), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n223), .B1(new_n220), .B2(new_n231), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n189), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G475), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(G475), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n217), .A2(KEYINPUT77), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n208), .A2(new_n211), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n195), .A2(new_n198), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n216), .A2(KEYINPUT19), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT19), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n245), .A3(new_n201), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n223), .B1(new_n247), .B2(new_n231), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n237), .B1(new_n248), .B2(new_n232), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(new_n237), .C1(new_n248), .C2(new_n232), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n236), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n256), .A2(G952), .ZN(new_n257));
  NAND2_X1  g071(.A1(G234), .A2(G237), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(G902), .A3(G953), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT21), .B(G898), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G478), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n266), .A2(KEYINPUT15), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT74), .B(G217), .Z(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n188), .A3(new_n256), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G122), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G122), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G107), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT13), .ZN(new_n280));
  INV_X1    g094(.A(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G143), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(G143), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G143), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G128), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n280), .ZN(new_n287));
  OAI21_X1  g101(.A(G134), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G134), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n286), .A2(new_n283), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n290), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n273), .A2(KEYINPUT14), .A3(G122), .ZN(new_n295));
  OAI211_X1 g109(.A(G107), .B(new_n295), .C1(new_n275), .C2(KEYINPUT14), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n278), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n270), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(new_n297), .A3(new_n270), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n267), .B1(new_n301), .B2(new_n189), .ZN(new_n302));
  INV_X1    g116(.A(new_n300), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n189), .B(new_n267), .C1(new_n303), .C2(new_n298), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n255), .A2(new_n265), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT83), .B(G469), .Z(new_n308));
  XNOR2_X1  g122(.A(G110), .B(G140), .ZN(new_n309));
  INV_X1    g123(.A(G227), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(G953), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n309), .B(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n277), .A2(G104), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n222), .A2(G107), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT78), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(KEYINPUT78), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n277), .A2(G104), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n201), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n285), .A2(G146), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(G128), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n281), .B1(new_n325), .B2(KEYINPUT1), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(G101), .B1(new_n316), .B2(new_n313), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n324), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n324), .A2(new_n332), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT65), .B1(new_n201), .B2(G143), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n325), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n328), .B1(new_n337), .B2(new_n330), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n333), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n289), .A2(G137), .ZN(new_n340));
  INV_X1    g154(.A(G137), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT66), .B1(new_n341), .B2(G134), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT11), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n343), .C1(new_n289), .C2(G137), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G131), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n345), .B1(new_n289), .B2(G137), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n197), .A3(new_n346), .A4(new_n340), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n339), .A2(KEYINPUT12), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n352), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT12), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(KEYINPUT0), .A2(G128), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n329), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT64), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(KEYINPUT0), .B2(G128), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n357), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n360), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n359), .B1(new_n337), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n317), .A2(new_n323), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(G101), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(new_n324), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n315), .B1(new_n316), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n222), .A2(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n320), .B2(new_n322), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n366), .B(G101), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n367), .A2(KEYINPUT79), .A3(new_n366), .A4(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n336), .A2(new_n325), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n325), .A2(KEYINPUT1), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(G128), .ZN(new_n384));
  INV_X1    g198(.A(new_n328), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(KEYINPUT68), .B(new_n328), .C1(new_n337), .C2(new_n330), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n334), .A2(new_n386), .A3(KEYINPUT10), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n333), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n348), .A2(new_n391), .A3(new_n351), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n391), .B1(new_n348), .B2(new_n351), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n379), .A2(new_n388), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n369), .A2(new_n378), .B1(new_n389), .B2(new_n333), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n388), .A4(new_n394), .ZN(new_n399));
  AOI221_X4 g213(.A(new_n312), .B1(new_n353), .B2(new_n356), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n312), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n399), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n398), .A2(new_n388), .B1(new_n348), .B2(new_n351), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n189), .B(new_n308), .C1(new_n400), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n401), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n356), .A2(new_n353), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n403), .B1(new_n397), .B2(new_n399), .ZN(new_n411));
  OAI22_X1  g225(.A1(new_n408), .A2(new_n410), .B1(new_n411), .B2(new_n401), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n189), .A4(new_n308), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n401), .B1(new_n402), .B2(new_n409), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n312), .B1(new_n397), .B2(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n403), .B1(new_n419), .B2(KEYINPUT82), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G469), .B1(new_n421), .B2(G902), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n190), .B(new_n307), .C1(new_n415), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G122), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT67), .B(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G116), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n273), .A2(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT2), .B(G113), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n432), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n367), .A2(G101), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n378), .A2(new_n427), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n429), .A2(KEYINPUT5), .A3(new_n430), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(G113), .C1(KEYINPUT5), .C2(new_n429), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n334), .A3(new_n435), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n368), .A2(new_n324), .B1(new_n433), .B2(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n427), .B1(new_n444), .B2(new_n378), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n426), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n378), .A2(new_n436), .A3(new_n438), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT85), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n448), .A2(new_n425), .A3(new_n442), .A4(new_n439), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(new_n426), .C1(new_n443), .C2(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(new_n213), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n384), .B2(new_n385), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n365), .B2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n256), .A2(G224), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT86), .Z(new_n457));
  XOR2_X1   g271(.A(new_n455), .B(new_n457), .Z(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n455), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n435), .ZN(new_n463));
  XOR2_X1   g277(.A(new_n463), .B(new_n334), .Z(new_n464));
  XNOR2_X1  g278(.A(new_n425), .B(KEYINPUT8), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n466), .B2(new_n449), .ZN(new_n467));
  OAI21_X1  g281(.A(G210), .B1(G237), .B2(G902), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n459), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n424), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT87), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n459), .A2(new_n467), .ZN(new_n473));
  INV_X1    g287(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n424), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G472), .A2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n289), .A2(G137), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n341), .A2(G134), .ZN(new_n484));
  OAI21_X1  g298(.A(G131), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n351), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n386), .A2(new_n486), .A3(new_n387), .ZN(new_n487));
  INV_X1    g301(.A(new_n436), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n357), .A2(KEYINPUT64), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n357), .B2(new_n361), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n285), .B2(G146), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n285), .A2(G146), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n382), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n490), .A2(new_n494), .B1(new_n358), .B2(new_n329), .ZN(new_n495));
  INV_X1    g309(.A(new_n351), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n484), .B1(new_n349), .B2(KEYINPUT11), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n197), .B1(new_n497), .B2(new_n346), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n487), .A2(new_n488), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n351), .B(new_n485), .C1(new_n384), .C2(new_n385), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n436), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n501), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT71), .B1(new_n500), .B2(new_n501), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT26), .B(G101), .Z(new_n509));
  NAND2_X1  g323(.A1(new_n191), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT72), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n506), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n500), .A2(KEYINPUT71), .A3(new_n501), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT72), .ZN(new_n519));
  INV_X1    g333(.A(new_n513), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n504), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n499), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n436), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT69), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT69), .A4(new_n436), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n513), .A3(new_n500), .A4(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n529), .A2(new_n500), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(KEYINPUT31), .A3(new_n513), .A4(new_n528), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n482), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT73), .B1(new_n536), .B2(KEYINPUT32), .ZN(new_n537));
  INV_X1    g351(.A(G472), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n526), .A2(new_n527), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n529), .A2(new_n500), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n520), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n502), .A2(new_n507), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n513), .A3(new_n515), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n500), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n488), .B1(new_n487), .B2(new_n499), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT28), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n520), .A2(new_n544), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n548), .A2(new_n516), .A3(new_n517), .A4(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(new_n189), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n536), .B2(KEYINPUT32), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT73), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n514), .A2(new_n521), .B1(new_n532), .B2(new_n534), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n482), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n537), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G234), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n268), .B1(new_n559), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n428), .B2(G128), .ZN(new_n562));
  OR2_X1    g376(.A1(G119), .A2(G128), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n428), .B2(new_n281), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(new_n561), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  OAI22_X1  g380(.A1(new_n565), .A2(G110), .B1(new_n566), .B2(new_n564), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n567), .A2(new_n238), .A3(new_n241), .A4(new_n226), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n565), .A2(G110), .B1(new_n566), .B2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n212), .A2(new_n217), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n187), .A2(new_n559), .A3(G953), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n568), .B(new_n579), .C1(new_n572), .C2(new_n573), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n189), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n578), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n560), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n580), .ZN(new_n586));
  INV_X1    g400(.A(new_n560), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n586), .A2(G902), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n423), .A2(new_n480), .A3(new_n558), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  AOI21_X1  g405(.A(new_n190), .B1(new_n415), .B2(new_n422), .ZN(new_n592));
  OAI21_X1  g406(.A(G472), .B1(new_n556), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n536), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  INV_X1    g410(.A(new_n471), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n252), .A2(new_n254), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n235), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n301), .A2(new_n600), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n300), .A2(KEYINPUT90), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n300), .A2(KEYINPUT90), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n603), .A2(KEYINPUT33), .A3(new_n299), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n266), .A2(G902), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n602), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n301), .A2(new_n189), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n266), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n599), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n597), .A2(new_n265), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  OR2_X1    g431(.A1(new_n248), .A2(new_n232), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n250), .A3(new_n237), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n236), .B1(new_n619), .B2(new_n252), .ZN(new_n620));
  INV_X1    g434(.A(new_n306), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n264), .B(KEYINPUT91), .Z(new_n623));
  NAND2_X1  g437(.A1(new_n597), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n596), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT35), .B(G107), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n583), .A2(new_n584), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n587), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n574), .B1(KEYINPUT36), .B2(new_n577), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n587), .A2(G902), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n568), .B(new_n632), .C1(new_n572), .C2(new_n573), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n307), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n480), .A2(new_n592), .A3(new_n595), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  XOR2_X1   g456(.A(new_n259), .B(KEYINPUT93), .Z(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n262), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n620), .A2(new_n621), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT94), .Z(new_n649));
  NOR2_X1   g463(.A1(new_n638), .A2(new_n471), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n558), .A2(new_n592), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XOR2_X1   g466(.A(new_n646), .B(KEYINPUT39), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n592), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n477), .B(KEYINPUT38), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n520), .B1(new_n546), .B2(new_n547), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n530), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n538), .B1(new_n658), .B2(new_n189), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n536), .B2(KEYINPUT32), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n537), .A2(new_n660), .A3(new_n557), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n255), .A2(new_n306), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n424), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n637), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n656), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n655), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT95), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NAND2_X1  g484(.A1(new_n613), .A2(new_n647), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n558), .A2(new_n592), .A3(new_n650), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  AND2_X1   g488(.A1(new_n558), .A2(new_n589), .ZN(new_n675));
  INV_X1    g489(.A(new_n614), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n402), .A2(new_n404), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n312), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n419), .A2(new_n409), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G469), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT96), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n412), .A2(new_n189), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT96), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(G469), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT97), .ZN(new_n687));
  INV_X1    g501(.A(new_n190), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .A4(new_n415), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n680), .A2(KEYINPUT96), .A3(new_n681), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n684), .B1(new_n683), .B2(G469), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n415), .B(new_n688), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT97), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n675), .A2(new_n676), .A3(new_n689), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n624), .A2(new_n622), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n675), .A2(new_n697), .A3(new_n689), .A4(new_n693), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  AND2_X1   g513(.A1(new_n558), .A2(new_n639), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n597), .A3(new_n689), .A4(new_n693), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(new_n623), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n471), .A2(new_n703), .A3(new_n663), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n542), .A2(new_n548), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n520), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n535), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT98), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n481), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n532), .A2(new_n534), .B1(new_n520), .B2(new_n705), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT98), .B1(new_n710), .B2(new_n482), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n589), .A2(new_n593), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n693), .A2(new_n704), .A3(new_n689), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT99), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NAND4_X1  g529(.A1(new_n593), .A2(new_n709), .A3(new_n637), .A4(new_n711), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n671), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n693), .A2(new_n717), .A3(new_n597), .A4(new_n689), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  AOI21_X1  g533(.A(new_n413), .B1(new_n680), .B2(new_n308), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n406), .A2(KEYINPUT84), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n422), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT100), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n190), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n477), .A2(KEYINPUT101), .A3(new_n664), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n469), .A2(new_n470), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n424), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n415), .A2(KEYINPUT100), .A3(new_n422), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n724), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n558), .A2(new_n589), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n734));
  INV_X1    g548(.A(new_n589), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n555), .B1(new_n556), .B2(new_n482), .ZN(new_n736));
  AOI211_X1 g550(.A(new_n735), .B(new_n671), .C1(new_n553), .C2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n729), .A3(new_n724), .A4(new_n730), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n733), .A2(new_n734), .B1(KEYINPUT42), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  INV_X1    g554(.A(new_n649), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n731), .A2(new_n732), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n289), .ZN(G36));
  NAND2_X1  g557(.A1(new_n611), .A2(new_n255), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT43), .Z(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n595), .A3(new_n638), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT44), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(KEYINPUT44), .ZN(new_n749));
  INV_X1    g563(.A(new_n729), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n421), .A2(KEYINPUT45), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT102), .ZN(new_n754));
  OAI21_X1  g568(.A(G469), .B1(new_n421), .B2(KEYINPUT45), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n681), .A2(new_n189), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT103), .B1(new_n758), .B2(KEYINPUT46), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT103), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n760), .B(new_n761), .C1(new_n756), .C2(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n759), .A2(new_n415), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n688), .ZN(new_n765));
  INV_X1    g579(.A(new_n653), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT104), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n768), .A3(new_n688), .A4(new_n653), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n752), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n341), .ZN(G39));
  NOR4_X1   g585(.A1(new_n750), .A2(new_n558), .A3(new_n589), .A4(new_n671), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT47), .B1(new_n764), .B2(new_n688), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n688), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n214), .ZN(G42));
  NAND2_X1  g592(.A1(new_n745), .A2(new_n644), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT111), .Z(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n712), .A3(new_n729), .ZN(new_n781));
  INV_X1    g595(.A(new_n776), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n774), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n686), .A2(new_n190), .A3(new_n415), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n693), .A2(new_n689), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(new_n729), .ZN(new_n787));
  INV_X1    g601(.A(new_n716), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n780), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT113), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n661), .A2(new_n735), .A3(new_n259), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n599), .A2(new_n611), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n664), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT112), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n780), .A2(new_n712), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n656), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT50), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n797), .A2(new_n799), .A3(KEYINPUT50), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n794), .B(new_n795), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT110), .B1(new_n785), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  OAI211_X1 g619(.A(KEYINPUT110), .B(new_n805), .C1(new_n785), .C2(new_n802), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n735), .B1(new_n553), .B2(new_n736), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n787), .A2(new_n807), .A3(new_n780), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n792), .A2(new_n613), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n786), .A2(new_n597), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n810), .B(new_n257), .C1(new_n811), .C2(new_n798), .ZN(new_n812));
  XOR2_X1   g626(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n813));
  AOI211_X1 g627(.A(new_n809), .B(new_n812), .C1(new_n808), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n804), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n620), .A2(new_n306), .A3(new_n647), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n637), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n729), .A3(new_n558), .A4(new_n592), .ZN(new_n820));
  INV_X1    g634(.A(new_n717), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n731), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n742), .A2(new_n822), .ZN(new_n823));
  AOI221_X4 g637(.A(new_n306), .B1(G475), .B2(new_n234), .C1(new_n252), .C2(new_n254), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT106), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n824), .A2(new_n825), .B1(new_n599), .B2(new_n611), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT106), .B1(new_n599), .B2(new_n306), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n703), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n472), .A3(new_n479), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n589), .A3(new_n592), .A4(new_n595), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n590), .A3(new_n640), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n823), .A2(new_n739), .A3(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n714), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n718), .A2(new_n651), .A3(new_n673), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n415), .A2(KEYINPUT100), .A3(new_n422), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT100), .B1(new_n415), .B2(new_n422), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n838), .A2(new_n839), .A3(new_n190), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n629), .A2(new_n636), .A3(new_n647), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n841), .A2(new_n471), .A3(new_n663), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n661), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n840), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n722), .A2(new_n723), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n688), .A3(new_n730), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n661), .A2(new_n842), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT109), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n837), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n837), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n718), .A2(new_n651), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n836), .A2(KEYINPUT53), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n837), .A2(new_n850), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n837), .A2(new_n850), .A3(new_n851), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n742), .A2(new_n831), .A3(new_n822), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n714), .A3(new_n739), .A4(new_n834), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n858), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n862), .A2(new_n864), .A3(new_n858), .ZN(new_n868));
  INV_X1    g682(.A(new_n835), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT108), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n869), .A2(new_n870), .A3(new_n739), .A4(new_n863), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n860), .A2(new_n861), .A3(new_n856), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n864), .A2(KEYINPUT108), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n868), .B1(new_n875), .B2(new_n858), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n867), .B1(new_n876), .B2(new_n866), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n815), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  OR4_X1    g692(.A1(new_n735), .A2(new_n664), .A3(new_n190), .A4(new_n744), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n686), .A2(new_n415), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n656), .B(new_n879), .C1(new_n880), .C2(KEYINPUT49), .ZN(new_n881));
  INV_X1    g695(.A(new_n661), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n881), .B(new_n882), .C1(KEYINPUT49), .C2(new_n880), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n256), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n189), .B1(new_n857), .B2(new_n865), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n450), .A2(new_n452), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n458), .ZN(new_n891));
  XNOR2_X1  g705(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n891), .B(new_n892), .Z(new_n893));
  OAI21_X1  g707(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n889), .B2(new_n893), .ZN(G51));
  AOI21_X1  g709(.A(new_n866), .B1(new_n857), .B2(new_n865), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n867), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n757), .B(KEYINPUT57), .Z(new_n900));
  OAI21_X1  g714(.A(new_n412), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n756), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n886), .B1(new_n901), .B2(new_n902), .ZN(G54));
  AND3_X1   g717(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n887), .B1(new_n904), .B2(new_n618), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n618), .B2(new_n904), .ZN(G60));
  AND3_X1   g720(.A1(new_n602), .A2(new_n605), .A3(new_n606), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n266), .A2(new_n189), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n908), .B(new_n909), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n877), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n907), .A2(new_n911), .ZN(new_n913));
  INV_X1    g727(.A(new_n867), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n896), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n887), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT117), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n886), .B1(new_n898), .B2(new_n913), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n872), .B1(new_n870), .B2(new_n836), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n920), .B2(new_n874), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n921), .B2(new_n868), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n910), .B1(new_n922), .B2(new_n867), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n918), .B(new_n919), .C1(new_n923), .C2(new_n907), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n924), .ZN(G63));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n857), .A2(new_n865), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  NAND4_X1  g744(.A1(new_n927), .A2(new_n633), .A3(new_n630), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n887), .ZN(new_n932));
  INV_X1    g746(.A(new_n930), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n857), .B2(new_n865), .ZN(new_n934));
  INV_X1    g748(.A(new_n586), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n926), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n927), .A2(new_n930), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n586), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n934), .A2(KEYINPUT119), .A3(new_n935), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n887), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n938), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n939), .A3(new_n586), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT119), .B1(new_n934), .B2(new_n935), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n949), .A2(KEYINPUT120), .A3(new_n944), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n937), .B1(new_n946), .B2(new_n950), .ZN(G66));
  INV_X1    g765(.A(new_n263), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n256), .B1(new_n952), .B2(G224), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n835), .A2(new_n831), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(new_n256), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n890), .B1(G898), .B2(new_n256), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  NOR2_X1   g772(.A1(new_n770), .A2(new_n777), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n826), .A2(new_n827), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n729), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n961), .A2(new_n732), .A3(new_n654), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n669), .A2(new_n837), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n669), .A2(KEYINPUT62), .A3(new_n837), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n524), .A2(new_n525), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT121), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n243), .A2(new_n245), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n742), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n739), .A2(new_n975), .A3(new_n837), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n767), .A2(new_n769), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n807), .A2(new_n597), .A3(new_n662), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n959), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n645), .A2(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT123), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n972), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n974), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n310), .B2(new_n645), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n968), .B2(new_n955), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n539), .A2(new_n540), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT124), .Z(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(new_n520), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n959), .A2(new_n954), .A3(new_n979), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n989), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n520), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n990), .A2(new_n993), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n541), .A2(new_n530), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n989), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n921), .B2(new_n868), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n998), .A2(new_n887), .A3(new_n1002), .ZN(G57));
endmodule


