

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U324 ( .A(n474), .B(n473), .ZN(n538) );
  XNOR2_X1 U325 ( .A(n452), .B(n451), .ZN(n527) );
  XNOR2_X1 U326 ( .A(n450), .B(KEYINPUT105), .ZN(n451) );
  AND2_X1 U327 ( .A1(G230GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U328 ( .A(KEYINPUT99), .B(KEYINPUT25), .ZN(n378) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n384) );
  XNOR2_X1 U330 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n473) );
  INV_X1 U331 ( .A(KEYINPUT37), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n314), .B(n292), .ZN(n315) );
  INV_X1 U333 ( .A(KEYINPUT55), .ZN(n481) );
  XNOR2_X1 U334 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U335 ( .A(n316), .B(n315), .ZN(n322) );
  XNOR2_X1 U336 ( .A(n481), .B(KEYINPUT121), .ZN(n482) );
  XNOR2_X1 U337 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U339 ( .A(n408), .B(KEYINPUT66), .Z(n543) );
  XNOR2_X1 U340 ( .A(n491), .B(G183GAT), .ZN(n492) );
  XNOR2_X1 U341 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U342 ( .A(n493), .B(n492), .ZN(G1350GAT) );
  XNOR2_X1 U343 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(G1GAT), .B(G15GAT), .Z(n446) );
  XOR2_X1 U345 ( .A(G43GAT), .B(KEYINPUT8), .Z(n294) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n427) );
  XOR2_X1 U348 ( .A(n446), .B(n427), .Z(n296) );
  NAND2_X1 U349 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U351 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n298) );
  XNOR2_X1 U352 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U355 ( .A(G36GAT), .B(G50GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G141GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U358 ( .A(G169GAT), .B(G197GAT), .Z(n304) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G8GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n513) );
  XOR2_X1 U363 ( .A(G148GAT), .B(KEYINPUT70), .Z(n359) );
  XNOR2_X1 U364 ( .A(G120GAT), .B(n359), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n309), .B(KEYINPUT33), .ZN(n324) );
  XNOR2_X1 U366 ( .A(G85GAT), .B(G106GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n310), .B(G99GAT), .ZN(n428) );
  INV_X1 U368 ( .A(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U369 ( .A(n428), .B(n311), .ZN(n316) );
  XOR2_X1 U370 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n313) );
  XNOR2_X1 U371 ( .A(KEYINPUT32), .B(KEYINPUT71), .ZN(n312) );
  XNOR2_X1 U372 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U373 ( .A(G71GAT), .B(G78GAT), .Z(n318) );
  XNOR2_X1 U374 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n432) );
  XOR2_X1 U376 ( .A(G176GAT), .B(G204GAT), .Z(n320) );
  XNOR2_X1 U377 ( .A(G92GAT), .B(G64GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n348) );
  XNOR2_X1 U379 ( .A(n432), .B(n348), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n577) );
  NOR2_X1 U382 ( .A1(n513), .A2(n577), .ZN(n494) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n325), .B(G113GAT), .ZN(n326) );
  XOR2_X1 U385 ( .A(n326), .B(KEYINPUT80), .Z(n328) );
  XNOR2_X1 U386 ( .A(G127GAT), .B(G134GAT), .ZN(n327) );
  XNOR2_X1 U387 ( .A(n328), .B(n327), .ZN(n399) );
  XOR2_X1 U388 ( .A(KEYINPUT17), .B(G169GAT), .Z(n330) );
  XNOR2_X1 U389 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n329) );
  XNOR2_X1 U390 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U391 ( .A(KEYINPUT83), .B(n331), .Z(n351) );
  XNOR2_X1 U392 ( .A(n399), .B(n351), .ZN(n341) );
  XOR2_X1 U393 ( .A(G183GAT), .B(G71GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(G15GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U396 ( .A(G99GAT), .B(G43GAT), .Z(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U398 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n337) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n338) );
  NAND2_X1 U401 ( .A1(G227GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n485) );
  INV_X1 U403 ( .A(n485), .ZN(n540) );
  XOR2_X1 U404 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n345) );
  XNOR2_X1 U405 ( .A(G211GAT), .B(G197GAT), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n363) );
  XOR2_X1 U407 ( .A(G183GAT), .B(G8GAT), .Z(n434) );
  XOR2_X1 U408 ( .A(KEYINPUT93), .B(n434), .Z(n347) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U411 ( .A(n349), .B(n348), .Z(n353) );
  XNOR2_X1 U412 ( .A(G218GAT), .B(G36GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n350), .B(G190GAT), .ZN(n415) );
  XNOR2_X1 U414 ( .A(n415), .B(n351), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n363), .B(n354), .ZN(n532) );
  NAND2_X1 U417 ( .A1(n540), .A2(n532), .ZN(n356) );
  INV_X1 U418 ( .A(KEYINPUT98), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n377) );
  XOR2_X1 U420 ( .A(KEYINPUT87), .B(KEYINPUT88), .Z(n358) );
  XNOR2_X1 U421 ( .A(G78GAT), .B(G204GAT), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U423 ( .A(n360), .B(n359), .Z(n362) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(G218GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U426 ( .A(n364), .B(n363), .Z(n366) );
  XOR2_X1 U427 ( .A(G162GAT), .B(G50GAT), .Z(n414) );
  XOR2_X1 U428 ( .A(G155GAT), .B(G22GAT), .Z(n433) );
  XNOR2_X1 U429 ( .A(n414), .B(n433), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n376) );
  XOR2_X1 U431 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n368) );
  XNOR2_X1 U432 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n374) );
  XOR2_X1 U434 ( .A(G141GAT), .B(KEYINPUT2), .Z(n370) );
  XNOR2_X1 U435 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n392) );
  XOR2_X1 U437 ( .A(n392), .B(KEYINPUT24), .Z(n372) );
  NAND2_X1 U438 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U440 ( .A(n374), .B(n373), .Z(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n479) );
  NOR2_X1 U442 ( .A1(n377), .A2(n479), .ZN(n379) );
  NAND2_X1 U443 ( .A1(n479), .A2(n485), .ZN(n382) );
  XOR2_X1 U444 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n380) );
  XNOR2_X1 U445 ( .A(KEYINPUT96), .B(n380), .ZN(n381) );
  XOR2_X1 U446 ( .A(n382), .B(n381), .Z(n570) );
  XNOR2_X1 U447 ( .A(n532), .B(KEYINPUT27), .ZN(n406) );
  AND2_X1 U448 ( .A1(n570), .A2(n406), .ZN(n383) );
  NOR2_X1 U449 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n385), .B(KEYINPUT100), .ZN(n404) );
  XOR2_X1 U451 ( .A(G148GAT), .B(G1GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G155GAT), .B(G57GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n389) );
  XNOR2_X1 U455 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n403) );
  XOR2_X1 U458 ( .A(G85GAT), .B(n392), .Z(n394) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U460 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U461 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n396) );
  XNOR2_X1 U462 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U464 ( .A(n398), .B(n397), .Z(n401) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n530) );
  NOR2_X1 U468 ( .A1(n404), .A2(n530), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n405), .B(KEYINPUT101), .ZN(n412) );
  NAND2_X1 U470 ( .A1(n406), .A2(n530), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n407), .B(KEYINPUT94), .ZN(n539) );
  XOR2_X1 U472 ( .A(n479), .B(KEYINPUT28), .Z(n408) );
  OR2_X1 U473 ( .A1(n540), .A2(n543), .ZN(n409) );
  NOR2_X1 U474 ( .A1(n539), .A2(n409), .ZN(n410) );
  XNOR2_X1 U475 ( .A(KEYINPUT95), .B(n410), .ZN(n411) );
  NAND2_X1 U476 ( .A1(n412), .A2(n411), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n413), .B(KEYINPUT102), .ZN(n497) );
  XOR2_X1 U478 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U479 ( .A(G134GAT), .B(G92GAT), .ZN(n416) );
  XNOR2_X1 U480 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U481 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n419) );
  NAND2_X1 U482 ( .A1(G232GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U483 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U485 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n423) );
  XNOR2_X1 U486 ( .A(KEYINPUT75), .B(KEYINPUT9), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(n424), .B(KEYINPUT65), .Z(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n465) );
  XNOR2_X1 U492 ( .A(n465), .B(KEYINPUT104), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n431), .B(KEYINPUT36), .ZN(n459) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U496 ( .A(G64GAT), .B(KEYINPUT76), .Z(n437) );
  NAND2_X1 U497 ( .A1(G231GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n444) );
  XOR2_X1 U500 ( .A(KEYINPUT15), .B(G211GAT), .Z(n441) );
  XNOR2_X1 U501 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n442), .B(KEYINPUT78), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n445), .B(KEYINPUT77), .ZN(n448) );
  XOR2_X1 U506 ( .A(G127GAT), .B(n446), .Z(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n467) );
  INV_X1 U508 ( .A(n467), .ZN(n458) );
  NOR2_X1 U509 ( .A1(n459), .A2(n467), .ZN(n449) );
  NAND2_X1 U510 ( .A1(n497), .A2(n449), .ZN(n452) );
  NAND2_X1 U511 ( .A1(n494), .A2(n527), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT38), .B(n453), .Z(n511) );
  NAND2_X1 U513 ( .A1(n511), .A2(n540), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n455) );
  INV_X1 U515 ( .A(G43GAT), .ZN(n454) );
  NOR2_X1 U516 ( .A1(n459), .A2(n458), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT45), .B(n460), .Z(n461) );
  NOR2_X1 U518 ( .A1(n461), .A2(n577), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n462), .A2(n513), .ZN(n472) );
  XNOR2_X1 U520 ( .A(KEYINPUT41), .B(n577), .ZN(n486) );
  NOR2_X1 U521 ( .A1(n513), .A2(n486), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT112), .ZN(n547) );
  NOR2_X1 U526 ( .A1(n468), .A2(n547), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT120), .B(n532), .Z(n475) );
  NOR2_X1 U531 ( .A1(n538), .A2(n475), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT54), .B(n476), .Z(n477) );
  NOR2_X1 U533 ( .A1(n530), .A2(n477), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT64), .ZN(n571) );
  INV_X1 U535 ( .A(n571), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n483) );
  NOR2_X1 U537 ( .A1(n485), .A2(n484), .ZN(n567) );
  INV_X1 U538 ( .A(n486), .ZN(n556) );
  NAND2_X1 U539 ( .A1(n567), .A2(n556), .ZN(n490) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT122), .Z(n488) );
  XNOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n487) );
  XNOR2_X1 U542 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U543 ( .A(n490), .B(n489), .ZN(G1349GAT) );
  NAND2_X1 U544 ( .A1(n567), .A2(n547), .ZN(n493) );
  XOR2_X1 U545 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n491) );
  INV_X1 U546 ( .A(n494), .ZN(n499) );
  NAND2_X1 U547 ( .A1(n467), .A2(n465), .ZN(n495) );
  XNOR2_X1 U548 ( .A(n495), .B(KEYINPUT16), .ZN(n496) );
  XNOR2_X1 U549 ( .A(KEYINPUT79), .B(n496), .ZN(n498) );
  NAND2_X1 U550 ( .A1(n498), .A2(n497), .ZN(n514) );
  NOR2_X1 U551 ( .A1(n499), .A2(n514), .ZN(n506) );
  NAND2_X1 U552 ( .A1(n506), .A2(n530), .ZN(n500) );
  XNOR2_X1 U553 ( .A(n500), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n501), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n532), .A2(n506), .ZN(n502) );
  XNOR2_X1 U556 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U558 ( .A1(n506), .A2(n540), .ZN(n503) );
  XNOR2_X1 U559 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U560 ( .A(G15GAT), .B(n505), .Z(G1326GAT) );
  NAND2_X1 U561 ( .A1(n543), .A2(n506), .ZN(n507) );
  XNOR2_X1 U562 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n509) );
  NAND2_X1 U564 ( .A1(n530), .A2(n511), .ZN(n508) );
  XNOR2_X1 U565 ( .A(n509), .B(n508), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n511), .A2(n532), .ZN(n510) );
  XNOR2_X1 U567 ( .A(n510), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n543), .A2(n511), .ZN(n512) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n512), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n517) );
  INV_X1 U571 ( .A(n513), .ZN(n572) );
  NOR2_X1 U572 ( .A1(n486), .A2(n572), .ZN(n528) );
  INV_X1 U573 ( .A(n528), .ZN(n515) );
  NOR2_X1 U574 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n523), .A2(n530), .ZN(n516) );
  XNOR2_X1 U576 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n518), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n532), .A2(n523), .ZN(n519) );
  XNOR2_X1 U579 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n521) );
  NAND2_X1 U581 ( .A1(n523), .A2(n540), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U585 ( .A1(n523), .A2(n543), .ZN(n524) );
  XNOR2_X1 U586 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U589 ( .A(n529), .B(KEYINPUT111), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n535), .A2(n530), .ZN(n531) );
  XNOR2_X1 U591 ( .A(n531), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n532), .A2(n535), .ZN(n533) );
  XNOR2_X1 U593 ( .A(n533), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n540), .A2(n535), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n534), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n543), .A2(n535), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n553) );
  NAND2_X1 U600 ( .A1(n553), .A2(n540), .ZN(n541) );
  XNOR2_X1 U601 ( .A(KEYINPUT116), .B(n541), .ZN(n542) );
  NOR2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n550), .A2(n572), .ZN(n544) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U606 ( .A1(n550), .A2(n556), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n547), .A2(n550), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n548), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n549), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  INV_X1 U612 ( .A(n465), .ZN(n566) );
  NAND2_X1 U613 ( .A1(n550), .A2(n566), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n553), .A2(n570), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT117), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n572), .A2(n562), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n560) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n558) );
  NAND2_X1 U621 ( .A1(n562), .A2(n556), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n562), .A2(n467), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U627 ( .A1(n562), .A2(n566), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n572), .A2(n567), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n583) );
  INV_X1 U636 ( .A(n583), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n580), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U642 ( .A1(n580), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n467), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n459), .A2(n583), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

