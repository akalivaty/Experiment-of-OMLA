

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n545), .A2(n548), .ZN(n793) );
  BUF_X1 U553 ( .A(n738), .Z(n522) );
  XNOR2_X1 U554 ( .A(n522), .B(n732), .ZN(n735) );
  NAND2_X1 U555 ( .A1(G8), .A2(n523), .ZN(n766) );
  NOR2_X1 U556 ( .A1(n699), .A2(G651), .ZN(n694) );
  XNOR2_X1 U557 ( .A(n565), .B(n564), .ZN(n698) );
  NAND2_X1 U558 ( .A1(n601), .A2(n526), .ZN(n602) );
  NOR2_X2 U559 ( .A1(G2104), .A2(G2105), .ZN(n586) );
  XNOR2_X2 U560 ( .A(n602), .B(KEYINPUT89), .ZN(G164) );
  INV_X1 U561 ( .A(KEYINPUT17), .ZN(n585) );
  AND2_X1 U562 ( .A1(n798), .A2(n529), .ZN(n799) );
  AND2_X1 U563 ( .A1(n782), .A2(n777), .ZN(n776) );
  OR2_X1 U564 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U565 ( .A1(n753), .A2(G299), .ZN(n751) );
  OR2_X1 U566 ( .A1(n764), .A2(n768), .ZN(n769) );
  AND2_X1 U567 ( .A1(n742), .A2(n741), .ZN(n746) );
  XNOR2_X1 U568 ( .A(n731), .B(KEYINPUT64), .ZN(n738) );
  AND2_X1 U569 ( .A1(n597), .A2(n596), .ZN(n601) );
  XNOR2_X1 U570 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U571 ( .A(n586), .B(n585), .ZN(n598) );
  AND2_X2 U572 ( .A1(G2105), .A2(G2104), .ZN(n915) );
  INV_X1 U573 ( .A(G2104), .ZN(n587) );
  AND2_X1 U574 ( .A1(n587), .A2(G2105), .ZN(n521) );
  AND2_X1 U575 ( .A1(n587), .A2(G2105), .ZN(n593) );
  BUF_X1 U576 ( .A(n738), .Z(n524) );
  NOR2_X2 U577 ( .A1(n591), .A2(n590), .ZN(G160) );
  NOR2_X2 U578 ( .A1(G1966), .A2(n766), .ZN(n786) );
  XNOR2_X2 U579 ( .A(n781), .B(KEYINPUT32), .ZN(n789) );
  BUF_X2 U580 ( .A(n738), .Z(n523) );
  NAND2_X1 U581 ( .A1(n552), .A2(n556), .ZN(n550) );
  XNOR2_X1 U582 ( .A(n799), .B(KEYINPUT107), .ZN(n800) );
  XNOR2_X1 U583 ( .A(n754), .B(KEYINPUT28), .ZN(n533) );
  AND2_X1 U584 ( .A1(n528), .A2(n554), .ZN(n553) );
  NAND2_X1 U585 ( .A1(n555), .A2(KEYINPUT105), .ZN(n554) );
  INV_X1 U586 ( .A(n791), .ZN(n555) );
  AND2_X1 U587 ( .A1(n791), .A2(n557), .ZN(n556) );
  INV_X1 U588 ( .A(G2105), .ZN(n582) );
  NAND2_X1 U589 ( .A1(n542), .A2(n540), .ZN(n539) );
  NAND2_X1 U590 ( .A1(n541), .A2(n850), .ZN(n540) );
  OR2_X1 U591 ( .A1(n810), .A2(KEYINPUT109), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n532), .B(n531), .ZN(n530) );
  INV_X1 U593 ( .A(KEYINPUT29), .ZN(n531) );
  XNOR2_X1 U594 ( .A(n773), .B(KEYINPUT104), .ZN(n774) );
  NAND2_X1 U595 ( .A1(n547), .A2(n546), .ZN(n545) );
  AND2_X1 U596 ( .A1(n550), .A2(n553), .ZN(n546) );
  XNOR2_X1 U597 ( .A(G1981), .B(G305), .ZN(n969) );
  INV_X1 U598 ( .A(n849), .ZN(n541) );
  AND2_X1 U599 ( .A1(n849), .A2(KEYINPUT109), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n810), .A2(n544), .ZN(n542) );
  XNOR2_X1 U601 ( .A(n637), .B(n636), .ZN(n643) );
  NOR2_X2 U602 ( .A1(n699), .A2(n563), .ZN(n686) );
  XNOR2_X1 U603 ( .A(KEYINPUT76), .B(n655), .ZN(n957) );
  XOR2_X1 U604 ( .A(KEYINPUT0), .B(G543), .Z(n699) );
  NOR2_X1 U605 ( .A1(G543), .A2(G651), .ZN(n685) );
  INV_X1 U606 ( .A(KEYINPUT87), .ZN(n594) );
  NAND2_X1 U607 ( .A1(n593), .A2(G126), .ZN(n595) );
  NAND2_X1 U608 ( .A1(n535), .A2(n582), .ZN(n592) );
  AND2_X1 U609 ( .A1(G102), .A2(G2104), .ZN(n535) );
  NAND2_X1 U610 ( .A1(n527), .A2(n582), .ZN(n583) );
  NAND2_X1 U611 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U612 ( .A1(n786), .A2(n785), .ZN(n525) );
  AND2_X1 U613 ( .A1(n600), .A2(n599), .ZN(n526) );
  AND2_X1 U614 ( .A1(G2104), .A2(G101), .ZN(n527) );
  NOR2_X1 U615 ( .A1(n766), .A2(n792), .ZN(n528) );
  AND2_X1 U616 ( .A1(n582), .A2(G2104), .ZN(n618) );
  XOR2_X1 U617 ( .A(n797), .B(KEYINPUT106), .Z(n529) );
  INV_X1 U618 ( .A(KEYINPUT105), .ZN(n557) );
  NAND2_X1 U619 ( .A1(n530), .A2(n759), .ZN(n782) );
  NAND2_X1 U620 ( .A1(n534), .A2(n533), .ZN(n532) );
  XNOR2_X1 U621 ( .A(n752), .B(KEYINPUT102), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n538), .A2(n536), .ZN(n865) );
  OR2_X1 U623 ( .A1(n811), .A2(n537), .ZN(n536) );
  NOR2_X1 U624 ( .A1(n543), .A2(n539), .ZN(n538) );
  AND2_X1 U625 ( .A1(n811), .A2(n544), .ZN(n543) );
  NAND2_X1 U626 ( .A1(n789), .A2(n551), .ZN(n547) );
  NOR2_X1 U627 ( .A1(n789), .A2(n549), .ZN(n548) );
  INV_X1 U628 ( .A(n556), .ZN(n549) );
  AND2_X1 U629 ( .A1(n788), .A2(KEYINPUT105), .ZN(n551) );
  NAND2_X1 U630 ( .A1(n789), .A2(n788), .ZN(n801) );
  INV_X1 U631 ( .A(n788), .ZN(n552) );
  XNOR2_X1 U632 ( .A(n592), .B(KEYINPUT88), .ZN(n597) );
  XOR2_X1 U633 ( .A(n808), .B(KEYINPUT98), .Z(n558) );
  XOR2_X1 U634 ( .A(KEYINPUT23), .B(n583), .Z(n559) );
  AND2_X1 U635 ( .A1(n523), .A2(G1341), .ZN(n560) );
  INV_X1 U636 ( .A(KEYINPUT99), .ZN(n732) );
  INV_X1 U637 ( .A(KEYINPUT27), .ZN(n733) );
  INV_X1 U638 ( .A(KEYINPUT31), .ZN(n773) );
  NAND2_X1 U639 ( .A1(n809), .A2(n558), .ZN(n810) );
  NAND2_X1 U640 ( .A1(G114), .A2(n915), .ZN(n599) );
  INV_X1 U641 ( .A(KEYINPUT15), .ZN(n653) );
  INV_X1 U642 ( .A(KEYINPUT14), .ZN(n636) );
  INV_X1 U643 ( .A(KEYINPUT109), .ZN(n850) );
  INV_X1 U644 ( .A(KEYINPUT1), .ZN(n564) );
  XNOR2_X1 U645 ( .A(n611), .B(KEYINPUT70), .ZN(G301) );
  XOR2_X1 U646 ( .A(KEYINPUT83), .B(KEYINPUT2), .Z(n562) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(G651), .ZN(n563) );
  NAND2_X1 U648 ( .A1(G73), .A2(n686), .ZN(n561) );
  XNOR2_X1 U649 ( .A(n562), .B(n561), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n694), .A2(G48), .ZN(n567) );
  NOR2_X1 U651 ( .A1(n563), .A2(G543), .ZN(n565) );
  NAND2_X1 U652 ( .A1(G61), .A2(n698), .ZN(n566) );
  NAND2_X1 U653 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U654 ( .A1(n685), .A2(G86), .ZN(n568) );
  XOR2_X1 U655 ( .A(KEYINPUT82), .B(n568), .Z(n569) );
  NOR2_X1 U656 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n572), .A2(n571), .ZN(G305) );
  NAND2_X1 U658 ( .A1(G53), .A2(n694), .ZN(n573) );
  XNOR2_X1 U659 ( .A(n573), .B(KEYINPUT72), .ZN(n580) );
  NAND2_X1 U660 ( .A1(G78), .A2(n686), .ZN(n575) );
  NAND2_X1 U661 ( .A1(G65), .A2(n698), .ZN(n574) );
  NAND2_X1 U662 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U663 ( .A1(G91), .A2(n685), .ZN(n576) );
  XNOR2_X1 U664 ( .A(KEYINPUT71), .B(n576), .ZN(n577) );
  NOR2_X1 U665 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(G299) );
  NAND2_X1 U667 ( .A1(G113), .A2(n915), .ZN(n581) );
  XNOR2_X1 U668 ( .A(n581), .B(KEYINPUT66), .ZN(n584) );
  NAND2_X1 U669 ( .A1(n584), .A2(n559), .ZN(n591) );
  BUF_X2 U670 ( .A(n598), .Z(n612) );
  NAND2_X1 U671 ( .A1(G137), .A2(n612), .ZN(n589) );
  NAND2_X1 U672 ( .A1(G125), .A2(n521), .ZN(n588) );
  NAND2_X1 U673 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n598), .A2(G138), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n685), .A2(G90), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G77), .A2(n686), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT9), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n694), .A2(G52), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G64), .A2(n698), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U682 ( .A(KEYINPUT69), .B(n608), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n611) );
  AND2_X1 U684 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U685 ( .A1(G111), .A2(n915), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G135), .A2(n612), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n521), .A2(G123), .ZN(n615) );
  XOR2_X1 U689 ( .A(KEYINPUT18), .B(n615), .Z(n616) );
  NOR2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n618), .A2(G99), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n1040) );
  XNOR2_X1 U693 ( .A(G2096), .B(n1040), .ZN(n621) );
  OR2_X1 U694 ( .A1(G2100), .A2(n621), .ZN(G156) );
  INV_X1 U695 ( .A(G57), .ZN(G237) );
  INV_X1 U696 ( .A(G132), .ZN(G219) );
  INV_X1 U697 ( .A(G82), .ZN(G220) );
  NAND2_X1 U698 ( .A1(n694), .A2(G51), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G63), .A2(n698), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U701 ( .A(KEYINPUT6), .B(n624), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n685), .A2(G89), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT4), .ZN(n627) );
  NAND2_X1 U704 ( .A1(G76), .A2(n686), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT5), .B(n628), .ZN(n629) );
  XNOR2_X1 U707 ( .A(KEYINPUT77), .B(n629), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT7), .B(n632), .Z(G168) );
  XOR2_X1 U710 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U711 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n634) );
  NAND2_X1 U712 ( .A1(G7), .A2(G661), .ZN(n633) );
  XNOR2_X1 U713 ( .A(n634), .B(n633), .ZN(G223) );
  XOR2_X1 U714 ( .A(G223), .B(KEYINPUT74), .Z(n867) );
  NAND2_X1 U715 ( .A1(n867), .A2(G567), .ZN(n635) );
  XOR2_X1 U716 ( .A(KEYINPUT11), .B(n635), .Z(G234) );
  NAND2_X1 U717 ( .A1(n698), .A2(G56), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n685), .A2(G81), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(KEYINPUT12), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G68), .A2(n686), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT13), .B(n641), .Z(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n694), .A2(G43), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n973) );
  INV_X1 U726 ( .A(G860), .ZN(n661) );
  OR2_X1 U727 ( .A1(n973), .A2(n661), .ZN(G153) );
  NAND2_X1 U728 ( .A1(G66), .A2(n698), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G92), .A2(n685), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G54), .A2(n694), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G79), .A2(n686), .ZN(n648) );
  XNOR2_X1 U733 ( .A(KEYINPUT75), .B(n648), .ZN(n649) );
  NOR2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U737 ( .A1(n957), .A2(G868), .ZN(n657) );
  INV_X1 U738 ( .A(G868), .ZN(n703) );
  NOR2_X1 U739 ( .A1(G301), .A2(n703), .ZN(n656) );
  NOR2_X1 U740 ( .A1(n657), .A2(n656), .ZN(G284) );
  NOR2_X1 U741 ( .A1(G286), .A2(n703), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT78), .ZN(n660) );
  NOR2_X1 U743 ( .A1(G299), .A2(G868), .ZN(n659) );
  NOR2_X1 U744 ( .A1(n660), .A2(n659), .ZN(G297) );
  NAND2_X1 U745 ( .A1(n661), .A2(G559), .ZN(n662) );
  INV_X1 U746 ( .A(n957), .ZN(n929) );
  NAND2_X1 U747 ( .A1(n662), .A2(n929), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U749 ( .A1(G868), .A2(n973), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n929), .A2(G868), .ZN(n664) );
  NOR2_X1 U751 ( .A1(G559), .A2(n664), .ZN(n665) );
  NOR2_X1 U752 ( .A1(n666), .A2(n665), .ZN(G282) );
  NAND2_X1 U753 ( .A1(G559), .A2(n929), .ZN(n711) );
  XNOR2_X1 U754 ( .A(n973), .B(n711), .ZN(n667) );
  NOR2_X1 U755 ( .A1(n667), .A2(G860), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G55), .A2(n694), .ZN(n668) );
  XNOR2_X1 U757 ( .A(n668), .B(KEYINPUT80), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n686), .A2(G80), .ZN(n669) );
  XOR2_X1 U759 ( .A(KEYINPUT79), .B(n669), .Z(n670) );
  NAND2_X1 U760 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U761 ( .A1(n685), .A2(G93), .ZN(n673) );
  NAND2_X1 U762 ( .A1(G67), .A2(n698), .ZN(n672) );
  NAND2_X1 U763 ( .A1(n673), .A2(n672), .ZN(n674) );
  OR2_X1 U764 ( .A1(n675), .A2(n674), .ZN(n706) );
  XOR2_X1 U765 ( .A(n676), .B(n706), .Z(G145) );
  NAND2_X1 U766 ( .A1(n694), .A2(G50), .ZN(n677) );
  XNOR2_X1 U767 ( .A(n677), .B(KEYINPUT84), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G62), .A2(n698), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U770 ( .A(KEYINPUT85), .B(n680), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n686), .A2(G75), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n685), .A2(G88), .ZN(n681) );
  AND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n684), .A2(n683), .ZN(G303) );
  INV_X1 U775 ( .A(G303), .ZN(G166) );
  NAND2_X1 U776 ( .A1(n685), .A2(G85), .ZN(n688) );
  NAND2_X1 U777 ( .A1(G72), .A2(n686), .ZN(n687) );
  NAND2_X1 U778 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U779 ( .A(KEYINPUT68), .B(n689), .Z(n693) );
  NAND2_X1 U780 ( .A1(n698), .A2(G60), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n694), .A2(G47), .ZN(n690) );
  AND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(G290) );
  NAND2_X1 U784 ( .A1(G49), .A2(n694), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G74), .A2(G651), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G87), .A2(n699), .ZN(n700) );
  XOR2_X1 U789 ( .A(KEYINPUT81), .B(n700), .Z(n701) );
  NAND2_X1 U790 ( .A1(n702), .A2(n701), .ZN(G288) );
  NAND2_X1 U791 ( .A1(n703), .A2(n706), .ZN(n714) );
  XNOR2_X1 U792 ( .A(G166), .B(G290), .ZN(n704) );
  XNOR2_X1 U793 ( .A(n704), .B(n973), .ZN(n705) );
  XOR2_X1 U794 ( .A(n706), .B(n705), .Z(n708) );
  XNOR2_X1 U795 ( .A(G288), .B(KEYINPUT19), .ZN(n707) );
  XNOR2_X1 U796 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U797 ( .A(n709), .B(G305), .Z(n710) );
  XNOR2_X1 U798 ( .A(G299), .B(n710), .ZN(n930) );
  XNOR2_X1 U799 ( .A(n930), .B(n711), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n712), .A2(G868), .ZN(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U802 ( .A(n715), .B(KEYINPUT86), .ZN(G295) );
  NAND2_X1 U803 ( .A1(G2084), .A2(G2078), .ZN(n716) );
  XOR2_X1 U804 ( .A(KEYINPUT20), .B(n716), .Z(n717) );
  NAND2_X1 U805 ( .A1(G2090), .A2(n717), .ZN(n718) );
  XNOR2_X1 U806 ( .A(KEYINPUT21), .B(n718), .ZN(n719) );
  NAND2_X1 U807 ( .A1(n719), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U808 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U809 ( .A1(G220), .A2(G219), .ZN(n720) );
  XOR2_X1 U810 ( .A(KEYINPUT22), .B(n720), .Z(n721) );
  NOR2_X1 U811 ( .A1(G218), .A2(n721), .ZN(n722) );
  NAND2_X1 U812 ( .A1(G96), .A2(n722), .ZN(n871) );
  NAND2_X1 U813 ( .A1(n871), .A2(G2106), .ZN(n726) );
  NAND2_X1 U814 ( .A1(G69), .A2(G120), .ZN(n723) );
  NOR2_X1 U815 ( .A1(G237), .A2(n723), .ZN(n724) );
  NAND2_X1 U816 ( .A1(G108), .A2(n724), .ZN(n872) );
  NAND2_X1 U817 ( .A1(n872), .A2(G567), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n873) );
  NAND2_X1 U819 ( .A1(G661), .A2(G483), .ZN(n727) );
  NOR2_X1 U820 ( .A1(n873), .A2(n727), .ZN(n870) );
  NAND2_X1 U821 ( .A1(n870), .A2(G36), .ZN(G176) );
  INV_X1 U822 ( .A(G301), .ZN(G171) );
  NOR2_X2 U823 ( .A1(G164), .A2(G1384), .ZN(n812) );
  NAND2_X1 U824 ( .A1(G160), .A2(G40), .ZN(n813) );
  INV_X1 U825 ( .A(n813), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n812), .A2(n730), .ZN(n731) );
  INV_X1 U827 ( .A(n735), .ZN(n755) );
  NAND2_X1 U828 ( .A1(G2072), .A2(n755), .ZN(n734) );
  XNOR2_X1 U829 ( .A(n734), .B(n733), .ZN(n737) );
  XOR2_X1 U830 ( .A(G1956), .B(KEYINPUT101), .Z(n984) );
  NAND2_X1 U831 ( .A1(n735), .A2(n984), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n753) );
  INV_X1 U833 ( .A(n524), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n739), .A2(G1996), .ZN(n740) );
  XNOR2_X1 U835 ( .A(n740), .B(KEYINPUT26), .ZN(n742) );
  NOR2_X1 U836 ( .A1(n560), .A2(n973), .ZN(n741) );
  NAND2_X1 U837 ( .A1(G2067), .A2(n755), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n523), .A2(G1348), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n747), .A2(n957), .ZN(n745) );
  NAND2_X1 U841 ( .A1(n746), .A2(n745), .ZN(n749) );
  OR2_X1 U842 ( .A1(n957), .A2(n747), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U844 ( .A1(G299), .A2(n753), .ZN(n754) );
  XNOR2_X1 U845 ( .A(KEYINPUT25), .B(G2078), .ZN(n1003) );
  NAND2_X1 U846 ( .A1(n1003), .A2(n755), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT100), .ZN(n758) );
  INV_X1 U848 ( .A(G1961), .ZN(n988) );
  NAND2_X1 U849 ( .A1(n523), .A2(n988), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n765), .A2(G171), .ZN(n759) );
  INV_X1 U852 ( .A(G8), .ZN(n764) );
  NOR2_X1 U853 ( .A1(G1971), .A2(n766), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n524), .A2(G2090), .ZN(n760) );
  NOR2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n762), .A2(G303), .ZN(n763) );
  OR2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n777) );
  NOR2_X1 U858 ( .A1(G171), .A2(n765), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n524), .A2(G2084), .ZN(n784) );
  NOR2_X1 U860 ( .A1(n786), .A2(n784), .ZN(n767) );
  XNOR2_X1 U861 ( .A(KEYINPUT103), .B(n767), .ZN(n768) );
  XNOR2_X1 U862 ( .A(n769), .B(KEYINPUT30), .ZN(n770) );
  NOR2_X1 U863 ( .A1(G168), .A2(n770), .ZN(n771) );
  NOR2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n775), .B(n774), .ZN(n783) );
  NAND2_X1 U866 ( .A1(n776), .A2(n783), .ZN(n780) );
  INV_X1 U867 ( .A(n777), .ZN(n778) );
  OR2_X1 U868 ( .A1(n778), .A2(G286), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n787) );
  AND2_X1 U871 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n787), .A2(n525), .ZN(n788) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n953) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n790) );
  NOR2_X1 U875 ( .A1(n953), .A2(n790), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n954) );
  INV_X1 U877 ( .A(n954), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n793), .B(KEYINPUT65), .ZN(n795) );
  INV_X1 U879 ( .A(KEYINPUT33), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U881 ( .A1(KEYINPUT33), .A2(n953), .ZN(n796) );
  NOR2_X1 U882 ( .A1(n766), .A2(n796), .ZN(n797) );
  NOR2_X1 U883 ( .A1(n800), .A2(n969), .ZN(n811) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G8), .A2(n802), .ZN(n803) );
  NAND2_X1 U886 ( .A1(n801), .A2(n803), .ZN(n804) );
  XNOR2_X1 U887 ( .A(n804), .B(KEYINPUT108), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n805), .A2(n766), .ZN(n809) );
  NOR2_X1 U889 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U890 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  NOR2_X1 U891 ( .A1(n766), .A2(n807), .ZN(n808) );
  NOR2_X1 U892 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U893 ( .A(n814), .B(KEYINPUT90), .ZN(n863) );
  INV_X1 U894 ( .A(n863), .ZN(n815) );
  XOR2_X1 U895 ( .A(G1986), .B(G290), .Z(n961) );
  OR2_X1 U896 ( .A1(n815), .A2(n961), .ZN(n848) );
  XNOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .ZN(n860) );
  NAND2_X1 U898 ( .A1(n618), .A2(G104), .ZN(n816) );
  XOR2_X1 U899 ( .A(KEYINPUT91), .B(n816), .Z(n818) );
  NAND2_X1 U900 ( .A1(n612), .A2(G140), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n819), .ZN(n825) );
  NAND2_X1 U903 ( .A1(n521), .A2(G128), .ZN(n820) );
  XNOR2_X1 U904 ( .A(n820), .B(KEYINPUT92), .ZN(n822) );
  NAND2_X1 U905 ( .A1(G116), .A2(n915), .ZN(n821) );
  NAND2_X1 U906 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U907 ( .A(KEYINPUT35), .B(n823), .Z(n824) );
  NOR2_X1 U908 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n826), .ZN(n924) );
  NOR2_X1 U910 ( .A1(n860), .A2(n924), .ZN(n1044) );
  NAND2_X1 U911 ( .A1(n1044), .A2(n863), .ZN(n858) );
  NAND2_X1 U912 ( .A1(G105), .A2(n618), .ZN(n827) );
  XNOR2_X1 U913 ( .A(n827), .B(KEYINPUT38), .ZN(n834) );
  NAND2_X1 U914 ( .A1(G117), .A2(n915), .ZN(n829) );
  NAND2_X1 U915 ( .A1(G141), .A2(n612), .ZN(n828) );
  NAND2_X1 U916 ( .A1(n829), .A2(n828), .ZN(n832) );
  NAND2_X1 U917 ( .A1(n521), .A2(G129), .ZN(n830) );
  XOR2_X1 U918 ( .A(KEYINPUT96), .B(n830), .Z(n831) );
  NOR2_X1 U919 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U920 ( .A1(n834), .A2(n833), .ZN(n899) );
  NAND2_X1 U921 ( .A1(G1996), .A2(n899), .ZN(n845) );
  NAND2_X1 U922 ( .A1(G95), .A2(n618), .ZN(n836) );
  NAND2_X1 U923 ( .A1(G131), .A2(n612), .ZN(n835) );
  NAND2_X1 U924 ( .A1(n836), .A2(n835), .ZN(n842) );
  NAND2_X1 U925 ( .A1(n915), .A2(G107), .ZN(n837) );
  XOR2_X1 U926 ( .A(KEYINPUT93), .B(n837), .Z(n839) );
  NAND2_X1 U927 ( .A1(n521), .A2(G119), .ZN(n838) );
  NAND2_X1 U928 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U929 ( .A(KEYINPUT94), .B(n840), .ZN(n841) );
  NOR2_X1 U930 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U931 ( .A(n843), .B(KEYINPUT95), .ZN(n927) );
  NAND2_X1 U932 ( .A1(G1991), .A2(n927), .ZN(n844) );
  NAND2_X1 U933 ( .A1(n845), .A2(n844), .ZN(n1045) );
  NAND2_X1 U934 ( .A1(n863), .A2(n1045), .ZN(n852) );
  NAND2_X1 U935 ( .A1(n858), .A2(n852), .ZN(n846) );
  XNOR2_X1 U936 ( .A(n846), .B(KEYINPUT97), .ZN(n847) );
  AND2_X1 U937 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U938 ( .A1(n899), .A2(G1996), .ZN(n851) );
  XNOR2_X1 U939 ( .A(n851), .B(KEYINPUT110), .ZN(n1035) );
  INV_X1 U940 ( .A(n852), .ZN(n855) );
  NOR2_X1 U941 ( .A1(G1991), .A2(n927), .ZN(n1043) );
  NOR2_X1 U942 ( .A1(G1986), .A2(G290), .ZN(n853) );
  NOR2_X1 U943 ( .A1(n1043), .A2(n853), .ZN(n854) );
  NOR2_X1 U944 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U945 ( .A1(n1035), .A2(n856), .ZN(n857) );
  XNOR2_X1 U946 ( .A(n857), .B(KEYINPUT39), .ZN(n859) );
  NAND2_X1 U947 ( .A1(n859), .A2(n858), .ZN(n861) );
  NAND2_X1 U948 ( .A1(n860), .A2(n924), .ZN(n1049) );
  NAND2_X1 U949 ( .A1(n861), .A2(n1049), .ZN(n862) );
  NAND2_X1 U950 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U951 ( .A(n866), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U952 ( .A1(G2106), .A2(n867), .ZN(G217) );
  AND2_X1 U953 ( .A1(G15), .A2(G2), .ZN(n868) );
  NAND2_X1 U954 ( .A1(G661), .A2(n868), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n869) );
  NAND2_X1 U956 ( .A1(n870), .A2(n869), .ZN(G188) );
  INV_X1 U958 ( .A(G120), .ZN(G236) );
  INV_X1 U959 ( .A(G96), .ZN(G221) );
  INV_X1 U960 ( .A(G69), .ZN(G235) );
  NOR2_X1 U961 ( .A1(n872), .A2(n871), .ZN(G325) );
  INV_X1 U962 ( .A(G325), .ZN(G261) );
  INV_X1 U963 ( .A(n873), .ZN(G319) );
  XOR2_X1 U964 ( .A(G2100), .B(G2096), .Z(n875) );
  XNOR2_X1 U965 ( .A(KEYINPUT42), .B(G2678), .ZN(n874) );
  XNOR2_X1 U966 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U967 ( .A(KEYINPUT43), .B(G2090), .Z(n877) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2072), .ZN(n876) );
  XNOR2_X1 U969 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U970 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U971 ( .A(G2084), .B(G2078), .ZN(n880) );
  XNOR2_X1 U972 ( .A(n881), .B(n880), .ZN(G227) );
  XOR2_X1 U973 ( .A(G1971), .B(G1966), .Z(n883) );
  XNOR2_X1 U974 ( .A(G1996), .B(G1981), .ZN(n882) );
  XNOR2_X1 U975 ( .A(n883), .B(n882), .ZN(n887) );
  XOR2_X1 U976 ( .A(G1956), .B(G1961), .Z(n885) );
  XNOR2_X1 U977 ( .A(G1986), .B(G1976), .ZN(n884) );
  XNOR2_X1 U978 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U979 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U980 ( .A(KEYINPUT113), .B(G2474), .ZN(n888) );
  XNOR2_X1 U981 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U982 ( .A(G1991), .B(KEYINPUT41), .Z(n890) );
  XNOR2_X1 U983 ( .A(n891), .B(n890), .ZN(G229) );
  NAND2_X1 U984 ( .A1(G124), .A2(n521), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n892), .B(KEYINPUT44), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n915), .A2(G112), .ZN(n893) );
  NAND2_X1 U987 ( .A1(n894), .A2(n893), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G100), .A2(n618), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G136), .A2(n612), .ZN(n895) );
  NAND2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U991 ( .A1(n898), .A2(n897), .ZN(G162) );
  XNOR2_X1 U992 ( .A(G162), .B(n899), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n900), .B(n1040), .ZN(n901) );
  XOR2_X1 U994 ( .A(n901), .B(KEYINPUT48), .Z(n903) );
  XNOR2_X1 U995 ( .A(G160), .B(KEYINPUT46), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n912) );
  NAND2_X1 U997 ( .A1(G118), .A2(n915), .ZN(n905) );
  NAND2_X1 U998 ( .A1(G130), .A2(n521), .ZN(n904) );
  NAND2_X1 U999 ( .A1(n905), .A2(n904), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(G106), .A2(n618), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n612), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1003 ( .A(KEYINPUT45), .B(n908), .Z(n909) );
  NOR2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1005 ( .A(n912), .B(n911), .Z(n923) );
  NAND2_X1 U1006 ( .A1(G103), .A2(n618), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n612), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n921) );
  NAND2_X1 U1009 ( .A1(n915), .A2(G115), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(n916), .B(KEYINPUT114), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(G127), .A2(n521), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1013 ( .A(KEYINPUT47), .B(n919), .Z(n920) );
  NOR2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n1030) );
  XNOR2_X1 U1015 ( .A(G164), .B(n1030), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(n923), .B(n922), .ZN(n925) );
  XOR2_X1 U1017 ( .A(n925), .B(n924), .Z(n926) );
  XNOR2_X1 U1018 ( .A(n927), .B(n926), .ZN(n928) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n928), .ZN(G395) );
  XNOR2_X1 U1020 ( .A(G286), .B(n929), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(n931), .B(n930), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(n932), .B(G301), .ZN(n933) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n933), .ZN(G397) );
  XNOR2_X1 U1024 ( .A(G2454), .B(G2427), .ZN(n943) );
  XOR2_X1 U1025 ( .A(KEYINPUT112), .B(G2430), .Z(n935) );
  XNOR2_X1 U1026 ( .A(G2443), .B(G2451), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(n935), .B(n934), .ZN(n939) );
  XOR2_X1 U1028 ( .A(G2446), .B(KEYINPUT111), .Z(n937) );
  XNOR2_X1 U1029 ( .A(G1348), .B(G1341), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(n937), .B(n936), .ZN(n938) );
  XOR2_X1 U1031 ( .A(n939), .B(n938), .Z(n941) );
  XNOR2_X1 U1032 ( .A(G2435), .B(G2438), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(n941), .B(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n943), .B(n942), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(G14), .ZN(n950) );
  NAND2_X1 U1036 ( .A1(G319), .A2(n950), .ZN(n947) );
  NOR2_X1 U1037 ( .A1(G227), .A2(G229), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT49), .B(n945), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n949) );
  NOR2_X1 U1040 ( .A1(G395), .A2(G397), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(G225) );
  INV_X1 U1042 ( .A(G225), .ZN(G308) );
  INV_X1 U1043 ( .A(G108), .ZN(G238) );
  INV_X1 U1044 ( .A(n950), .ZN(G401) );
  XOR2_X1 U1045 ( .A(KEYINPUT56), .B(G16), .Z(n978) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G166), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT122), .ZN(n966) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G299), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n964) );
  XNOR2_X1 U1051 ( .A(n988), .B(G301), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT120), .ZN(n959) );
  XOR2_X1 U1053 ( .A(n957), .B(G1348), .Z(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT123), .B(n967), .ZN(n972) );
  XOR2_X1 U1060 ( .A(G1966), .B(G168), .Z(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n970), .Z(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT124), .B(n976), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n1027) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n979), .B(G4), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(G1981), .B(G6), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G1341), .B(G19), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(G20), .B(n984), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n987), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(n988), .B(G5), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n1000) );
  XOR2_X1 U1079 ( .A(G1966), .B(G21), .Z(n998) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1976), .B(G23), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n996), .B(KEYINPUT58), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n1001), .Z(n1002) );
  NOR2_X1 U1090 ( .A1(G16), .A2(n1002), .ZN(n1024) );
  XOR2_X1 U1091 ( .A(G1996), .B(G32), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1003), .B(G27), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(KEYINPUT119), .B(n1006), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(G1991), .B(G25), .Z(n1007) );
  NAND2_X1 U1096 ( .A1(G28), .A2(n1007), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT118), .B(G2072), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(G33), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G26), .B(G2067), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1015), .Z(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT54), .B(G34), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G2084), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G35), .B(G2090), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(KEYINPUT55), .B(n1021), .Z(n1022) );
  NOR2_X1 U1110 ( .A1(G29), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(G11), .A2(n1025), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1114 ( .A(n1028), .B(KEYINPUT126), .ZN(n1058) );
  XNOR2_X1 U1115 ( .A(G164), .B(G2078), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(n1029), .B(KEYINPUT117), .ZN(n1032) );
  XOR2_X1 U1117 ( .A(G2072), .B(n1030), .Z(n1031) );
  NOR2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT50), .B(n1033), .ZN(n1039) );
  XOR2_X1 U1120 ( .A(G2090), .B(G162), .Z(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1122 ( .A(KEYINPUT116), .B(n1036), .Z(n1037) );
  XNOR2_X1 U1123 ( .A(KEYINPUT51), .B(n1037), .ZN(n1038) );
  NAND2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1052) );
  XNOR2_X1 U1125 ( .A(G160), .B(G2084), .ZN(n1041) );
  NAND2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NOR2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1047) );
  NOR2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1129 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1130 ( .A(KEYINPUT115), .B(n1048), .ZN(n1050) );
  NAND2_X1 U1131 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NOR2_X1 U1132 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  XNOR2_X1 U1133 ( .A(KEYINPUT52), .B(n1053), .ZN(n1055) );
  INV_X1 U1134 ( .A(KEYINPUT55), .ZN(n1054) );
  NAND2_X1 U1135 ( .A1(n1055), .A2(n1054), .ZN(n1056) );
  NAND2_X1 U1136 ( .A1(n1056), .A2(G29), .ZN(n1057) );
  NAND2_X1 U1137 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XOR2_X1 U1138 ( .A(KEYINPUT62), .B(n1059), .Z(G311) );
  INV_X1 U1139 ( .A(G311), .ZN(G150) );
endmodule

