//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  AND3_X1   g003(.A1(new_n203), .A2(KEYINPUT73), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT73), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(new_n203), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n208), .A3(new_n203), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n214), .B(new_n202), .C1(new_n205), .C2(new_n206), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n217));
  NAND2_X1  g016(.A1(G226gat), .A2(G233gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT26), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n220), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT27), .B(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT28), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT28), .B(new_n230), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n228), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n234), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n222), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT23), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G176gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n219), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n227), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n244), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n257), .A2(new_n260), .A3(new_n227), .A4(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n238), .A2(new_n243), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n217), .B(new_n218), .C1(new_n263), .C2(KEYINPUT29), .ZN(new_n264));
  AND4_X1   g063(.A1(new_n227), .A2(new_n257), .A3(new_n260), .A4(new_n261), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT65), .B(G176gat), .Z(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT64), .B(G169gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT23), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(new_n227), .A3(new_n257), .A4(new_n247), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n265), .B1(new_n269), .B2(new_n244), .ZN(new_n270));
  INV_X1    g069(.A(new_n236), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT76), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n218), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n259), .A2(new_n262), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT76), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n236), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n242), .B2(new_n228), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n217), .B1(new_n283), .B2(new_n218), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n216), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n272), .A2(new_n282), .A3(new_n218), .A4(new_n276), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n273), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n213), .A2(new_n215), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n294), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(KEYINPUT30), .A3(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n285), .A2(new_n290), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G141gat), .ZN(new_n304));
  INV_X1    g103(.A(G141gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G148gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT2), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(KEYINPUT77), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G155gat), .B(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n304), .B2(new_n306), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n312), .B1(new_n316), .B2(new_n310), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(new_n313), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n312), .A3(new_n310), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n325));
  OAI21_X1  g124(.A(G113gat), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G113gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G120gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(KEYINPUT70), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G134gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G127gat), .ZN(new_n331));
  INV_X1    g130(.A(G127gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n328), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT67), .B1(new_n332), .B2(G134gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n330), .A3(G127gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n340), .A2(new_n342), .A3(new_n333), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G113gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT1), .B1(new_n328), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n339), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n340), .A2(new_n342), .A3(new_n333), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(KEYINPUT68), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n329), .A2(new_n338), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT4), .B1(new_n323), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n350), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n314), .A2(new_n317), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n337), .ZN(new_n355));
  INV_X1    g154(.A(new_n335), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n329), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n354), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n353), .A2(new_n354), .A3(new_n357), .A4(KEYINPUT78), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT5), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n359), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT4), .B1(new_n361), .B2(new_n362), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n354), .A3(new_n357), .A4(KEYINPUT4), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n369), .B(new_n364), .C1(new_n351), .C2(new_n323), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT5), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(new_n362), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n373));
  INV_X1    g172(.A(new_n354), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n364), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n367), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378));
  INV_X1    g177(.A(G85gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  INV_X1    g183(.A(new_n382), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n367), .C1(new_n371), .C2(new_n376), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n302), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n289), .B1(new_n282), .B2(new_n322), .ZN(new_n396));
  INV_X1    g195(.A(new_n212), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n207), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n212), .B(new_n202), .C1(new_n206), .C2(new_n205), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n282), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n354), .B1(new_n320), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n395), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n213), .B2(new_n215), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n374), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n404));
  INV_X1    g203(.A(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n322), .A2(new_n282), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n216), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G22gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n402), .B2(new_n408), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n394), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n402), .A2(new_n408), .A3(KEYINPUT80), .A4(new_n409), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n410), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n416), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n413), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n422), .A2(KEYINPUT82), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(KEYINPUT82), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n390), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n281), .A2(new_n373), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n238), .A2(new_n243), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n351), .A3(new_n274), .ZN(new_n428));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT72), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n426), .B2(new_n428), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT34), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n429), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n281), .A2(new_n373), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n351), .B1(new_n427), .B2(new_n274), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT34), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT32), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n432), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n434), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n434), .B2(new_n440), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n431), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n443), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n438), .B2(new_n444), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n439), .B1(new_n438), .B2(KEYINPUT32), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT34), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n431), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n440), .A3(new_n446), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT36), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n383), .A2(KEYINPUT83), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n377), .A2(new_n462), .A3(new_n382), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n364), .B1(new_n359), .B2(new_n363), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n372), .A2(new_n364), .A3(new_n375), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT39), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n382), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n470), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n464), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n302), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT84), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n464), .A2(new_n473), .A3(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n478), .A2(new_n302), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n422), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n386), .A2(new_n384), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n388), .A2(KEYINPUT85), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n296), .B1(new_n299), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n288), .B2(new_n216), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n289), .B1(new_n278), .B2(new_n284), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT38), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n297), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT38), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n291), .A2(KEYINPUT37), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n482), .B1(new_n487), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n460), .B1(new_n481), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n486), .A3(new_n485), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n416), .A2(new_n418), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n413), .A2(new_n506), .B1(new_n449), .B2(new_n457), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(new_n302), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n298), .A2(new_n301), .B1(new_n387), .B2(new_n388), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n510), .B(new_n511), .C1(new_n507), .C2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n302), .A2(new_n458), .A3(new_n389), .A4(new_n422), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT87), .B1(new_n514), .B2(KEYINPUT35), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  OR2_X1    g324(.A1(G57gat), .A2(G64gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G57gat), .A2(G64gat), .ZN(new_n527));
  AND2_X1   g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(KEYINPUT9), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n528), .ZN(new_n531));
  NOR2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n535), .B(new_n529), .C1(new_n530), .C2(new_n528), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(KEYINPUT93), .A3(new_n536), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n525), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(new_n332), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n543), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT96), .B(G155gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n541), .A2(new_n542), .ZN(new_n553));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n551), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n551), .B2(new_n552), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n566), .A2(KEYINPUT88), .A3(KEYINPUT15), .ZN(new_n567));
  OR3_X1    g366(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n568), .A2(new_n569), .B1(G29gat), .B2(G36gat), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT15), .B1(new_n566), .B2(KEYINPUT88), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT89), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n574), .A2(new_n575), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT17), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n379), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G99gat), .B(G106gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT98), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n578), .A2(new_n592), .A3(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G134gat), .B(G162gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n577), .A2(new_n588), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n596), .B1(new_n594), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n565), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n564), .A3(new_n598), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n560), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n578), .A2(new_n525), .ZN(new_n606));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT91), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n525), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n577), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(new_n577), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n608), .B(KEYINPUT13), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n606), .A2(KEYINPUT18), .A3(new_n609), .A4(new_n611), .ZN(new_n617));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618));
  INV_X1    g417(.A(G197gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT11), .B(G169gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n616), .B2(new_n617), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n588), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n539), .A2(new_n627), .A3(new_n540), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n588), .A2(new_n537), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n541), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT100), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n636), .B1(new_n628), .B2(new_n630), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n637), .A2(new_n641), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n541), .A2(new_n632), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n635), .B1(new_n647), .B2(new_n631), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n640), .B1(new_n648), .B2(new_n642), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n626), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n605), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n517), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n389), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g456(.A1(new_n654), .A2(new_n476), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n658), .B2(new_n518), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g460(.A(KEYINPUT42), .B(new_n659), .S(new_n661), .Z(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n654), .B2(new_n458), .ZN(new_n663));
  INV_X1    g462(.A(new_n459), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT102), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n654), .B2(new_n666), .ZN(G1326gat));
  OR2_X1    g466(.A1(new_n423), .A2(new_n424), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n654), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  AOI21_X1  g470(.A(new_n604), .B1(new_n501), .B2(new_n516), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n560), .A2(new_n652), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G29gat), .A3(new_n389), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n516), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n509), .B(new_n679), .C1(new_n513), .C2(new_n515), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n500), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(new_n604), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n672), .A2(KEYINPUT44), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n673), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n389), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n676), .A2(new_n686), .ZN(G1328gat));
  NOR3_X1   g486(.A1(new_n674), .A2(G36gat), .A3(new_n302), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT46), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n685), .B2(new_n302), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1329gat));
  INV_X1    g490(.A(new_n458), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n674), .A2(G43gat), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n684), .A2(new_n664), .A3(new_n673), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G43gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g495(.A(G50gat), .B1(new_n685), .B2(new_n422), .ZN(new_n697));
  INV_X1    g496(.A(new_n668), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n674), .A2(G50gat), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(KEYINPUT48), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n697), .A2(KEYINPUT104), .A3(KEYINPUT48), .A4(new_n699), .ZN(new_n703));
  OAI21_X1  g502(.A(G50gat), .B1(new_n685), .B2(new_n698), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(new_n699), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n702), .B(new_n703), .C1(KEYINPUT48), .C2(new_n705), .ZN(G1331gat));
  NOR4_X1   g505(.A1(new_n681), .A2(new_n626), .A3(new_n651), .A4(new_n605), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n655), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g508(.A1(new_n707), .A2(new_n476), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(G1333gat));
  NAND2_X1  g513(.A1(new_n707), .A2(new_n664), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n458), .B(KEYINPUT105), .Z(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(G71gat), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n715), .A2(G71gat), .B1(new_n707), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n707), .A2(new_n668), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n560), .A2(new_n626), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n651), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n682), .A2(new_n683), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT106), .A4(new_n724), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(new_n379), .A3(new_n389), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n678), .A2(new_n680), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n501), .ZN(new_n732));
  INV_X1    g531(.A(new_n604), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n722), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n733), .A4(new_n722), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n681), .A2(new_n604), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(KEYINPUT107), .A3(KEYINPUT51), .A4(new_n722), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n737), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n745), .A2(new_n655), .A3(new_n650), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n730), .B1(new_n746), .B2(new_n379), .ZN(G1336gat));
  NOR2_X1   g546(.A1(new_n302), .A2(G92gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n650), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n681), .A2(new_n604), .A3(new_n723), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n750), .B2(KEYINPUT51), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n752), .A3(new_n735), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n749), .B1(new_n754), .B2(new_n743), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n302), .B1(new_n727), .B2(new_n728), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n755), .A2(KEYINPUT110), .B1(new_n756), .B2(new_n584), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n758), .B(new_n749), .C1(new_n754), .C2(new_n743), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n650), .A3(new_n748), .ZN(new_n761));
  XNOR2_X1  g560(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n684), .A2(new_n476), .A3(new_n724), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(G92gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(new_n765), .ZN(G1337gat));
  XOR2_X1   g565(.A(KEYINPUT112), .B(G99gat), .Z(new_n767));
  NOR2_X1   g566(.A1(new_n692), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n745), .A2(new_n650), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n729), .B2(new_n459), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  OR3_X1    g570(.A1(new_n422), .A2(new_n651), .A3(G106gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n745), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n725), .A2(new_n775), .A3(new_n422), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n725), .B2(new_n422), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  OAI21_X1  g579(.A(G106gat), .B1(new_n729), .B2(new_n698), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n754), .A2(new_n743), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n782), .B2(new_n773), .ZN(new_n783));
  AOI22_X1  g582(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n783), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n624), .A2(new_n625), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n560), .A2(new_n785), .A3(new_n651), .A4(new_n604), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n609), .B1(new_n606), .B2(new_n611), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n614), .A2(new_n615), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n622), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND4_X1   g589(.A1(new_n787), .A2(new_n601), .A3(new_n603), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n646), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n633), .B2(new_n636), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n647), .A2(new_n631), .A3(KEYINPUT114), .A4(new_n635), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT54), .A4(new_n637), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n641), .B1(new_n648), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n792), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n796), .A2(new_n798), .A3(new_n802), .A4(KEYINPUT55), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n796), .A2(new_n798), .A3(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n650), .A3(new_n790), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n785), .B2(new_n806), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n791), .A2(new_n807), .B1(new_n809), .B2(new_n604), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n786), .B1(new_n810), .B2(new_n560), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n655), .A3(new_n507), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT116), .Z(new_n813));
  NAND4_X1  g612(.A1(new_n813), .A2(new_n327), .A3(new_n302), .A4(new_n626), .ZN(new_n814));
  INV_X1    g613(.A(new_n811), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n668), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n476), .A2(new_n389), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n816), .A2(new_n458), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n785), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT117), .Z(G1340gat));
  OR2_X1    g620(.A1(new_n324), .A2(new_n325), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n813), .A2(new_n822), .A3(new_n302), .A4(new_n650), .ZN(new_n823));
  OAI21_X1  g622(.A(G120gat), .B1(new_n818), .B2(new_n651), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT118), .ZN(G1341gat));
  INV_X1    g625(.A(new_n560), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n818), .A2(new_n332), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT119), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n302), .A3(new_n560), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n332), .ZN(G1342gat));
  AND4_X1   g630(.A1(new_n330), .A2(new_n813), .A3(new_n302), .A4(new_n733), .ZN(new_n832));
  XOR2_X1   g631(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n818), .B2(new_n604), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n791), .A2(new_n807), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n806), .A2(KEYINPUT121), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n801), .A2(new_n805), .A3(new_n841), .A4(new_n803), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n626), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n808), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n733), .B1(new_n844), .B2(KEYINPUT122), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n846), .A3(new_n808), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n786), .B1(new_n848), .B2(new_n560), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n668), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n811), .A2(new_n482), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(KEYINPUT57), .ZN(new_n853));
  INV_X1    g652(.A(new_n817), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n664), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n851), .A2(new_n626), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n852), .A2(new_n856), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n305), .A3(new_n626), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n859), .B(new_n863), .C1(new_n860), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n862), .A2(new_n303), .A3(new_n650), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n849), .B2(new_n668), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n852), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n811), .A2(KEYINPUT124), .A3(KEYINPUT57), .A4(new_n482), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n650), .B(new_n855), .C1(new_n871), .C2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n303), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n850), .A2(new_n873), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(KEYINPUT125), .A3(new_n650), .A4(new_n855), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n870), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n853), .B(new_n856), .C1(new_n850), .C2(KEYINPUT57), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT59), .B(new_n303), .C1(new_n885), .C2(new_n650), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n869), .B1(new_n884), .B2(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(G155gat), .B1(new_n862), .B2(new_n560), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n827), .A2(new_n308), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n885), .B2(new_n889), .ZN(G1346gat));
  NAND3_X1  g689(.A1(new_n733), .A2(new_n302), .A3(new_n459), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G162gat), .A3(new_n422), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n811), .A2(new_n655), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n885), .A2(new_n733), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n309), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n476), .A2(new_n389), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n716), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n816), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G169gat), .B1(new_n898), .B2(new_n785), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n507), .A2(new_n476), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(KEYINPUT126), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(KEYINPUT126), .ZN(new_n902));
  NOR4_X1   g701(.A1(new_n815), .A2(new_n655), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n267), .A3(new_n626), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n904), .ZN(G1348gat));
  NOR3_X1   g704(.A1(new_n898), .A2(new_n266), .A3(new_n651), .ZN(new_n906));
  AOI21_X1  g705(.A(G176gat), .B1(new_n903), .B2(new_n650), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(G183gat), .B1(new_n898), .B2(new_n827), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n903), .A2(new_n229), .A3(new_n560), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n816), .A2(new_n733), .A3(new_n897), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G190gat), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n230), .A3(new_n733), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n664), .A2(new_n896), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n852), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n619), .A3(new_n626), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n880), .B2(new_n881), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(new_n626), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(new_n619), .ZN(G1352gat));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n924), .A2(new_n929), .A3(new_n650), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT62), .Z(new_n931));
  AOI211_X1 g730(.A(new_n651), .B(new_n923), .C1(new_n880), .C2(new_n881), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n929), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n209), .A3(new_n560), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n926), .A2(new_n560), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n924), .B2(new_n733), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n604), .A2(new_n210), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n926), .B2(new_n940), .ZN(G1355gat));
endmodule


