

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599;

  NOR2_X2 U326 ( .A1(n543), .A2(n542), .ZN(n557) );
  INV_X1 U327 ( .A(n546), .ZN(n368) );
  XOR2_X1 U328 ( .A(n315), .B(n314), .Z(n572) );
  OR2_X1 U329 ( .A1(n542), .A2(n369), .ZN(n294) );
  XNOR2_X1 U330 ( .A(KEYINPUT116), .B(KEYINPUT45), .ZN(n470) );
  XNOR2_X1 U331 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G106GAT), .ZN(n407) );
  NAND2_X1 U333 ( .A1(n368), .A2(n490), .ZN(n369) );
  XNOR2_X1 U334 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U335 ( .A(n419), .B(n418), .ZN(n422) );
  XNOR2_X1 U336 ( .A(n401), .B(KEYINPUT105), .ZN(n429) );
  INV_X1 U337 ( .A(KEYINPUT96), .ZN(n323) );
  XOR2_X1 U338 ( .A(G176GAT), .B(G64GAT), .Z(n449) );
  XNOR2_X1 U339 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U340 ( .A(n326), .B(n325), .ZN(n331) );
  NOR2_X1 U341 ( .A1(n531), .A2(n498), .ZN(n465) );
  NOR2_X1 U342 ( .A1(n574), .A2(n490), .ZN(n579) );
  XNOR2_X1 U343 ( .A(n465), .B(KEYINPUT38), .ZN(n515) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n491) );
  XNOR2_X1 U345 ( .A(n466), .B(G43GAT), .ZN(n467) );
  XNOR2_X1 U346 ( .A(n492), .B(n491), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n468), .B(n467), .ZN(G1330GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT83), .B(KEYINPUT0), .Z(n296) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT82), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n342) );
  XOR2_X1 U351 ( .A(n342), .B(G190GAT), .Z(n298) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n299), .B(G99GAT), .Z(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n301) );
  XNOR2_X1 U356 ( .A(KEYINPUT85), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(KEYINPUT18), .B(n302), .Z(n319) );
  XOR2_X1 U359 ( .A(G71GAT), .B(G120GAT), .Z(n304) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n319), .B(n305), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n315) );
  XOR2_X1 U364 ( .A(G176GAT), .B(KEYINPUT87), .Z(n309) );
  XNOR2_X1 U365 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U367 ( .A(KEYINPUT20), .B(G127GAT), .Z(n311) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U370 ( .A(n313), .B(n312), .Z(n314) );
  XOR2_X1 U371 ( .A(n449), .B(G92GAT), .Z(n317) );
  XOR2_X1 U372 ( .A(G169GAT), .B(G8GAT), .Z(n436) );
  XNOR2_X1 U373 ( .A(n436), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(n319), .B(n318), .Z(n321) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n326) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n322), .B(G218GAT), .ZN(n413) );
  XNOR2_X1 U380 ( .A(n413), .B(KEYINPUT76), .ZN(n324) );
  XNOR2_X1 U381 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n327), .B(KEYINPUT21), .ZN(n328) );
  XOR2_X1 U383 ( .A(n328), .B(KEYINPUT90), .Z(n330) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(G211GAT), .ZN(n329) );
  XOR2_X1 U385 ( .A(n330), .B(n329), .Z(n364) );
  XOR2_X1 U386 ( .A(n331), .B(n364), .Z(n332) );
  XNOR2_X1 U387 ( .A(n332), .B(KEYINPUT27), .ZN(n374) );
  XOR2_X1 U388 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n334) );
  XNOR2_X1 U389 ( .A(G162GAT), .B(G85GAT), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U391 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n336) );
  XNOR2_X1 U392 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U394 ( .A(n338), .B(n337), .Z(n347) );
  XOR2_X1 U395 ( .A(KEYINPUT3), .B(KEYINPUT91), .Z(n340) );
  XNOR2_X1 U396 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(G141GAT), .B(n341), .Z(n363) );
  XOR2_X1 U399 ( .A(KEYINPUT4), .B(n342), .Z(n344) );
  NAND2_X1 U400 ( .A1(G225GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n363), .B(n345), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U404 ( .A(G1GAT), .B(G127GAT), .Z(n393) );
  XOR2_X1 U405 ( .A(n348), .B(n393), .Z(n351) );
  XNOR2_X1 U406 ( .A(G29GAT), .B(G134GAT), .ZN(n402) );
  XNOR2_X1 U407 ( .A(G120GAT), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n349), .B(G57GAT), .ZN(n458) );
  XOR2_X1 U409 ( .A(n402), .B(n458), .Z(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n378) );
  XNOR2_X1 U411 ( .A(KEYINPUT95), .B(n378), .ZN(n534) );
  NAND2_X1 U412 ( .A1(n374), .A2(n534), .ZN(n542) );
  XOR2_X1 U413 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n353) );
  XNOR2_X1 U414 ( .A(G218GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(n354), .B(G148GAT), .Z(n356) );
  XOR2_X1 U417 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U418 ( .A(G22GAT), .B(n423), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U420 ( .A(G78GAT), .B(G204GAT), .Z(n358) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n459) );
  XOR2_X1 U423 ( .A(KEYINPUT23), .B(n459), .Z(n360) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U426 ( .A(n362), .B(n361), .Z(n366) );
  XOR2_X1 U427 ( .A(n364), .B(n363), .Z(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n486) );
  XNOR2_X1 U429 ( .A(n486), .B(KEYINPUT64), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n367), .B(KEYINPUT28), .ZN(n546) );
  INV_X1 U431 ( .A(n572), .ZN(n490) );
  XOR2_X1 U432 ( .A(KEYINPUT97), .B(n294), .Z(n380) );
  XNOR2_X1 U433 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n372) );
  INV_X1 U434 ( .A(n332), .ZN(n484) );
  NOR2_X1 U435 ( .A1(n484), .A2(n490), .ZN(n370) );
  NOR2_X1 U436 ( .A1(n486), .A2(n370), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n376) );
  NAND2_X1 U438 ( .A1(n490), .A2(n486), .ZN(n373) );
  XOR2_X1 U439 ( .A(n373), .B(KEYINPUT26), .Z(n584) );
  NAND2_X1 U440 ( .A1(n374), .A2(n584), .ZN(n375) );
  NAND2_X1 U441 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U442 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U443 ( .A1(n380), .A2(n379), .ZN(n495) );
  XOR2_X1 U444 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n382) );
  XNOR2_X1 U445 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U447 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n384) );
  XNOR2_X1 U448 ( .A(KEYINPUT77), .B(KEYINPUT79), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n400) );
  XOR2_X1 U451 ( .A(G78GAT), .B(G155GAT), .Z(n388) );
  XNOR2_X1 U452 ( .A(G183GAT), .B(G211GAT), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U454 ( .A(KEYINPUT76), .B(G64GAT), .Z(n390) );
  XNOR2_X1 U455 ( .A(G8GAT), .B(G57GAT), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U457 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U458 ( .A(G15GAT), .B(G22GAT), .Z(n435) );
  XOR2_X1 U459 ( .A(G71GAT), .B(KEYINPUT13), .Z(n450) );
  XOR2_X1 U460 ( .A(n450), .B(n393), .Z(n395) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n435), .B(n396), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n400), .B(n399), .Z(n593) );
  INV_X1 U466 ( .A(n593), .ZN(n493) );
  NAND2_X1 U467 ( .A1(n495), .A2(n493), .ZN(n401) );
  INV_X1 U468 ( .A(n402), .ZN(n427) );
  INV_X1 U469 ( .A(G85GAT), .ZN(n403) );
  NAND2_X1 U470 ( .A1(G92GAT), .A2(n403), .ZN(n406) );
  INV_X1 U471 ( .A(G92GAT), .ZN(n404) );
  NAND2_X1 U472 ( .A1(n404), .A2(G85GAT), .ZN(n405) );
  NAND2_X1 U473 ( .A1(n406), .A2(n405), .ZN(n408) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n451) );
  INV_X1 U475 ( .A(KEYINPUT73), .ZN(n409) );
  XNOR2_X1 U476 ( .A(n451), .B(n409), .ZN(n411) );
  NAND2_X1 U477 ( .A1(G232GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n419) );
  XNOR2_X1 U479 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n412), .B(KEYINPUT7), .ZN(n444) );
  XNOR2_X1 U481 ( .A(n444), .B(n413), .ZN(n417) );
  XOR2_X1 U482 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n415) );
  XNOR2_X1 U483 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n414) );
  XOR2_X1 U484 ( .A(n415), .B(n414), .Z(n416) );
  INV_X1 U485 ( .A(n422), .ZN(n421) );
  INV_X1 U486 ( .A(n423), .ZN(n420) );
  NAND2_X1 U487 ( .A1(n421), .A2(n420), .ZN(n425) );
  NAND2_X1 U488 ( .A1(n423), .A2(n422), .ZN(n424) );
  NAND2_X1 U489 ( .A1(n425), .A2(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(n427), .B(n426), .Z(n476) );
  INV_X1 U491 ( .A(KEYINPUT75), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n476), .B(n428), .ZN(n553) );
  XNOR2_X1 U493 ( .A(KEYINPUT36), .B(n553), .ZN(n469) );
  BUF_X1 U494 ( .A(n469), .Z(n595) );
  NAND2_X1 U495 ( .A1(n429), .A2(n595), .ZN(n430) );
  XOR2_X1 U496 ( .A(KEYINPUT37), .B(n430), .Z(n531) );
  XOR2_X1 U497 ( .A(G141GAT), .B(G197GAT), .Z(n432) );
  XNOR2_X1 U498 ( .A(G29GAT), .B(G113GAT), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT66), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U501 ( .A(KEYINPUT65), .B(KEYINPUT30), .ZN(n433) );
  XNOR2_X1 U502 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U503 ( .A(G50GAT), .B(G36GAT), .Z(n438) );
  XNOR2_X1 U504 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U506 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U507 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U508 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U509 ( .A(n443), .B(KEYINPUT67), .Z(n446) );
  XNOR2_X1 U510 ( .A(n444), .B(KEYINPUT29), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U512 ( .A(n448), .B(n447), .Z(n517) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n463) );
  XOR2_X1 U514 ( .A(n451), .B(KEYINPUT68), .Z(n453) );
  NAND2_X1 U515 ( .A1(G230GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U517 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n455) );
  XNOR2_X1 U518 ( .A(KEYINPUT32), .B(KEYINPUT69), .ZN(n454) );
  XNOR2_X1 U519 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U520 ( .A(n457), .B(n456), .Z(n461) );
  XNOR2_X1 U521 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U523 ( .A(n463), .B(n462), .Z(n589) );
  OR2_X1 U524 ( .A1(n517), .A2(n589), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n464), .B(KEYINPUT72), .ZN(n498) );
  NAND2_X1 U526 ( .A1(n572), .A2(n515), .ZN(n468) );
  XOR2_X1 U527 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n466) );
  NAND2_X1 U528 ( .A1(n593), .A2(n469), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n589), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT117), .ZN(n474) );
  INV_X1 U531 ( .A(n517), .ZN(n585) );
  NOR2_X1 U532 ( .A1(n474), .A2(n585), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n475), .B(KEYINPUT118), .ZN(n482) );
  XOR2_X1 U534 ( .A(KEYINPUT41), .B(n589), .Z(n561) );
  NAND2_X1 U535 ( .A1(n585), .A2(n561), .ZN(n477) );
  XNOR2_X1 U536 ( .A(KEYINPUT46), .B(n477), .ZN(n478) );
  NAND2_X1 U537 ( .A1(n478), .A2(n493), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n476), .A2(n479), .ZN(n480) );
  XOR2_X1 U539 ( .A(KEYINPUT47), .B(n480), .Z(n481) );
  NOR2_X1 U540 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(KEYINPUT48), .ZN(n543) );
  NOR2_X1 U542 ( .A1(n484), .A2(n543), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT54), .B(n485), .ZN(n582) );
  INV_X1 U544 ( .A(n534), .ZN(n581) );
  INV_X1 U545 ( .A(n486), .ZN(n487) );
  AND2_X1 U546 ( .A1(n581), .A2(n487), .ZN(n488) );
  AND2_X1 U547 ( .A1(n582), .A2(n488), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT55), .ZN(n574) );
  NAND2_X1 U549 ( .A1(n579), .A2(n553), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n500) );
  NOR2_X1 U551 ( .A1(n493), .A2(n553), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(KEYINPUT16), .ZN(n496) );
  NAND2_X1 U553 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT99), .B(n497), .Z(n518) );
  NOR2_X1 U555 ( .A1(n498), .A2(n518), .ZN(n507) );
  NAND2_X1 U556 ( .A1(n507), .A2(n534), .ZN(n499) );
  XNOR2_X1 U557 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n501), .Z(G1324GAT) );
  XOR2_X1 U559 ( .A(G8GAT), .B(KEYINPUT101), .Z(n503) );
  NAND2_X1 U560 ( .A1(n507), .A2(n332), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U563 ( .A1(n507), .A2(n572), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  XOR2_X1 U566 ( .A(G22GAT), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U567 ( .A1(n507), .A2(n546), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1327GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n511) );
  NAND2_X1 U570 ( .A1(n515), .A2(n534), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G29GAT), .B(n512), .ZN(G1328GAT) );
  NAND2_X1 U573 ( .A1(n515), .A2(n332), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n513), .B(KEYINPUT106), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G36GAT), .B(n514), .ZN(G1329GAT) );
  NAND2_X1 U576 ( .A1(n515), .A2(n546), .ZN(n516) );
  XNOR2_X1 U577 ( .A(n516), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n521) );
  XNOR2_X1 U579 ( .A(KEYINPUT108), .B(n561), .ZN(n571) );
  NAND2_X1 U580 ( .A1(n517), .A2(n571), .ZN(n532) );
  NOR2_X1 U581 ( .A1(n532), .A2(n518), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT109), .B(n519), .Z(n526) );
  NAND2_X1 U583 ( .A1(n526), .A2(n534), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NAND2_X1 U586 ( .A1(n332), .A2(n526), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U588 ( .A(G71GAT), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n572), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n528) );
  NAND2_X1 U592 ( .A1(n526), .A2(n546), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n530) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT113), .Z(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1335GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT114), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n539), .A2(n534), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n539), .A2(n332), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U602 ( .A(G99GAT), .B(KEYINPUT115), .Z(n538) );
  NAND2_X1 U603 ( .A1(n572), .A2(n539), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n539), .A2(n546), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT44), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  NAND2_X1 U608 ( .A1(n572), .A2(n557), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(n544), .Z(n545) );
  NOR2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n585), .A2(n554), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n549) );
  NAND2_X1 U614 ( .A1(n554), .A2(n571), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G120GAT), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U617 ( .A1(n593), .A2(n554), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(KEYINPUT50), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n559) );
  AND2_X1 U624 ( .A1(n584), .A2(n557), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n567), .A2(n585), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U629 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n593), .A2(n567), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n476), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U637 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n579), .A2(n585), .ZN(n570) );
  XNOR2_X1 U639 ( .A(G169GAT), .B(n570), .ZN(G1348GAT) );
  XOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT125), .Z(n576) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n578) );
  XOR2_X1 U644 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(G1349GAT) );
  NAND2_X1 U646 ( .A1(n593), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n587) );
  AND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  AND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n596) );
  NAND2_X1 U651 ( .A1(n596), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G197GAT), .B(n588), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n591) );
  NAND2_X1 U655 ( .A1(n596), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(G204GAT), .B(n592), .ZN(G1353GAT) );
  NAND2_X1 U658 ( .A1(n593), .A2(n596), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n594), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U660 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n598) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U663 ( .A(G218GAT), .B(n599), .ZN(G1355GAT) );
endmodule

