//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G128), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT73), .B(G110), .Z(new_n194));
  INV_X1    g008(.A(KEYINPUT74), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n195), .B1(new_n193), .B2(new_n194), .ZN(new_n197));
  XNOR2_X1  g011(.A(G119), .B(G128), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  OAI211_X1 g013(.A(new_n196), .B(new_n197), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT71), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .A4(KEYINPUT16), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT71), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n202), .A2(new_n204), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n200), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT22), .B(G137), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n215), .B(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n212), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n193), .A2(G110), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n199), .A2(new_n198), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT72), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n226), .B(new_n223), .C1(new_n210), .C2(new_n219), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n214), .B(new_n218), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT76), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(KEYINPUT71), .C1(KEYINPUT16), .C2(new_n202), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n212), .B1(new_n231), .B2(new_n206), .ZN(new_n232));
  INV_X1    g046(.A(new_n219), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n224), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n226), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n220), .A2(KEYINPUT72), .A3(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT76), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n238), .A3(new_n214), .A4(new_n218), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n214), .B1(new_n225), .B2(new_n227), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT75), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n214), .C1(new_n225), .C2(new_n227), .ZN(new_n244));
  INV_X1    g058(.A(new_n218), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n240), .A2(new_n246), .A3(KEYINPUT25), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(G234), .B2(new_n247), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n240), .A2(new_n246), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(G902), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT77), .Z(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G237), .A2(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(KEYINPUT2), .A2(G113), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NOR3_X1   g085(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G116), .B(G119), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n274), .B(new_n269), .C1(new_n271), .C2(new_n272), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n212), .A2(G143), .ZN(new_n280));
  INV_X1    g094(.A(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  NOR2_X1   g098(.A1(KEYINPUT0), .A2(G128), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n288));
  XNOR2_X1  g102(.A(G143), .B(G146), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n284), .ZN(new_n290));
  AND4_X1   g104(.A1(new_n288), .A2(new_n280), .A3(new_n282), .A4(new_n284), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n293));
  INV_X1    g107(.A(G137), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT11), .B1(new_n294), .B2(G134), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(G134), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OR2_X1    g111(.A1(KEYINPUT66), .A2(G137), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT66), .A2(G137), .ZN(new_n299));
  AND2_X1   g113(.A1(KEYINPUT11), .A2(G134), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT67), .A2(G131), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT67), .A2(G131), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n297), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(KEYINPUT66), .A2(G137), .ZN(new_n306));
  NOR2_X1   g120(.A1(KEYINPUT66), .A2(G137), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n308), .A2(new_n300), .B1(new_n296), .B2(new_n295), .ZN(new_n309));
  INV_X1    g123(.A(G131), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT64), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n280), .A2(new_n282), .A3(new_n284), .A4(new_n288), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n287), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n293), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT1), .B1(new_n281), .B2(G146), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n283), .A2(G128), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n280), .B(new_n282), .C1(KEYINPUT1), .C2(new_n191), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G134), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n306), .B2(new_n307), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n310), .B1(new_n324), .B2(new_n296), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n305), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n279), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n313), .A2(new_n314), .B1(new_n283), .B2(new_n286), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n311), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n330), .A2(new_n327), .A3(new_n279), .ZN(new_n331));
  OAI211_X1 g145(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n328), .C2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n311), .B1(new_n329), .B2(new_n316), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n278), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n327), .A3(new_n279), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n333), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n268), .B(new_n332), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT70), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n331), .B1(new_n278), .B2(new_n336), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n341), .B(new_n340), .C1(new_n345), .C2(new_n333), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n268), .A4(new_n332), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n330), .A2(new_n327), .A3(KEYINPUT30), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n320), .A2(new_n321), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n297), .A2(new_n301), .A3(new_n304), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n351), .A2(new_n352), .A3(new_n325), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n297), .A2(new_n301), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G131), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n292), .A2(KEYINPUT65), .B1(new_n355), .B2(new_n305), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n356), .B2(new_n317), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n278), .B(new_n350), .C1(new_n357), .C2(KEYINPUT30), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n338), .A3(new_n267), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT31), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT31), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n338), .A4(new_n267), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G472), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n247), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n368), .A2(G472), .A3(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n330), .A2(new_n327), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n278), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n338), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT28), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT29), .A3(new_n267), .A4(new_n340), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(new_n247), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n268), .B1(new_n346), .B2(new_n332), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n330), .A2(new_n327), .A3(KEYINPUT30), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(new_n336), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n331), .B1(new_n381), .B2(new_n278), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n378), .B1(new_n382), .B2(new_n267), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n376), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n365), .A2(new_n370), .B1(G472), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n262), .B1(new_n369), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G214), .B1(G237), .B2(G902), .ZN(new_n387));
  XNOR2_X1  g201(.A(G110), .B(G122), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G101), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT3), .A3(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(G107), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n276), .A2(new_n277), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n394), .A2(KEYINPUT3), .A3(G104), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT3), .B1(new_n394), .B2(G104), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT79), .A3(G101), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n394), .A2(G104), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n393), .B2(new_n395), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n407), .B2(new_n390), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n399), .B1(new_n407), .B2(new_n390), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n404), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT80), .B1(new_n394), .B2(G104), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n392), .A3(G107), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n394), .A2(G104), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n188), .A2(G116), .ZN(new_n418));
  INV_X1    g232(.A(G116), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G119), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT5), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n419), .A2(G119), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n424), .A3(G113), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n390), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n417), .A2(new_n277), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT68), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT2), .ZN(new_n431));
  INV_X1    g245(.A(G113), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n270), .B1(KEYINPUT2), .B2(G113), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n422), .B2(new_n423), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n434), .A2(new_n274), .B1(new_n435), .B2(new_n421), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT84), .A3(new_n426), .A4(new_n417), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n389), .B1(new_n411), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n400), .A2(new_n410), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n440), .A2(new_n388), .A3(new_n429), .A4(new_n437), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G125), .B1(new_n320), .B2(new_n321), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n292), .B2(G125), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n216), .A2(G224), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(new_n389), .C1(new_n411), .C2(new_n438), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n442), .A2(new_n446), .A3(KEYINPUT85), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n445), .B1(KEYINPUT87), .B2(KEYINPUT7), .ZN(new_n456));
  AND2_X1   g270(.A1(KEYINPUT87), .A2(KEYINPUT7), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n203), .B1(new_n315), .B2(new_n287), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n455), .B(new_n459), .C1(new_n460), .C2(new_n443), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n277), .A2(new_n425), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n426), .A4(new_n417), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n417), .A2(new_n463), .A3(new_n426), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n436), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n388), .B(KEYINPUT8), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n461), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n292), .A2(G125), .ZN(new_n470));
  INV_X1    g284(.A(new_n443), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(KEYINPUT7), .A3(new_n471), .A4(new_n445), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT88), .B1(new_n444), .B2(new_n458), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n469), .A2(new_n441), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n454), .B1(new_n474), .B2(new_n247), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n473), .A2(new_n461), .A3(new_n468), .A4(new_n472), .ZN(new_n476));
  INV_X1    g290(.A(new_n441), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n454), .B(new_n247), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT90), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n453), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n453), .B2(new_n480), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n387), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT20), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n392), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n211), .B(new_n212), .ZN(new_n492));
  INV_X1    g306(.A(G237), .ZN(new_n493));
  AND4_X1   g307(.A1(G143), .A2(new_n493), .A3(new_n216), .A4(G214), .ZN(new_n494));
  AOI21_X1  g308(.A(G143), .B1(new_n263), .B2(G214), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(KEYINPUT18), .A2(G131), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n497), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT91), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n216), .A3(G214), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n281), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n263), .A2(G143), .A3(G214), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n500), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT92), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n509), .B(new_n500), .C1(new_n501), .C2(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n499), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n304), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n496), .A2(new_n304), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT17), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT67), .B(G131), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT17), .B(new_n517), .C1(new_n494), .C2(new_n495), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT94), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n512), .B2(KEYINPUT17), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n219), .B(new_n210), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n516), .B1(new_n522), .B2(KEYINPUT95), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n518), .B(KEYINPUT94), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n219), .A4(new_n210), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n491), .B(new_n511), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n508), .A2(new_n510), .ZN(new_n528));
  INV_X1    g342(.A(new_n499), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n211), .B(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n232), .B1(new_n212), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT93), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n515), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n490), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n487), .B(new_n488), .C1(new_n527), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n541));
  INV_X1    g355(.A(new_n516), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n526), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n490), .A3(new_n530), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n530), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n491), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n547), .A2(KEYINPUT96), .A3(new_n487), .A4(new_n488), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n511), .B1(new_n523), .B2(new_n526), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n537), .B1(new_n549), .B2(new_n490), .ZN(new_n550));
  INV_X1    g364(.A(new_n488), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT20), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n540), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n216), .A2(G952), .ZN(new_n554));
  NAND2_X1  g368(.A1(G234), .A2(G237), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(G902), .A3(G953), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(G128), .B(G143), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n323), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT98), .ZN(new_n565));
  XOR2_X1   g379(.A(G116), .B(G122), .Z(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G107), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(KEYINPUT13), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n281), .A2(G128), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(G134), .C1(KEYINPUT13), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT9), .B(G234), .Z(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT78), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n573), .A2(new_n253), .A3(G953), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n563), .B(new_n323), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n419), .A2(KEYINPUT14), .A3(G122), .ZN(new_n576));
  OAI211_X1 g390(.A(G107), .B(new_n576), .C1(new_n566), .C2(KEYINPUT14), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n577), .C1(G107), .C2(new_n566), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n571), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n574), .B1(new_n571), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n247), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI221_X1 g398(.A(new_n247), .B1(KEYINPUT15), .B2(new_n582), .C1(new_n579), .C2(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n490), .B1(new_n543), .B2(new_n530), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n247), .B1(new_n527), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT97), .B(G475), .Z(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n553), .A2(new_n562), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT82), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n417), .A2(new_n426), .A3(new_n321), .A4(new_n320), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n417), .A2(new_n426), .B1(new_n320), .B2(new_n321), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n311), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT12), .B1(new_n311), .B2(KEYINPUT81), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI221_X1 g413(.A(new_n311), .B1(KEYINPUT81), .B2(KEYINPUT12), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n398), .A2(new_n399), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n410), .A2(new_n329), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n310), .B1(new_n297), .B2(new_n301), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n352), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n322), .A2(KEYINPUT10), .A3(new_n426), .A4(new_n417), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n603), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(G110), .B(G140), .ZN(new_n611));
  INV_X1    g425(.A(G227), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(G953), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n410), .A2(new_n329), .A3(new_n602), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n608), .A2(new_n607), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n311), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n610), .A2(new_n614), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n593), .B(G469), .C1(new_n620), .C2(G902), .ZN(new_n621));
  INV_X1    g435(.A(G469), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT83), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n609), .A2(new_n623), .A3(new_n615), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n609), .B2(new_n615), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n417), .A2(new_n426), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n351), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n605), .B1(new_n627), .B2(new_n594), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n598), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n615), .B1(new_n619), .B2(new_n609), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n622), .B(new_n247), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n619), .A2(new_n615), .A3(new_n609), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n617), .A2(new_n618), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n634), .A2(new_n605), .B1(new_n599), .B2(new_n600), .ZN(new_n635));
  OAI211_X1 g449(.A(G469), .B(new_n633), .C1(new_n635), .C2(new_n615), .ZN(new_n636));
  NAND2_X1  g450(.A1(G469), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n636), .A2(KEYINPUT82), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n621), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G221), .B1(new_n573), .B2(G902), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n486), .A2(new_n592), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n386), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  INV_X1    g458(.A(new_n254), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n250), .B2(new_n251), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n641), .A2(new_n260), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n366), .B1(new_n365), .B2(new_n247), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n363), .B1(new_n344), .B2(new_n348), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n649), .A2(G472), .A3(G902), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n255), .A2(new_n261), .A3(new_n640), .A4(new_n639), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n649), .B2(G902), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n367), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT99), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT100), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n552), .A2(new_n548), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n551), .B1(new_n544), .B2(new_n546), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT96), .B1(new_n661), .B2(new_n487), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n591), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT101), .B(G478), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n581), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n579), .A2(new_n580), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT33), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n582), .A2(G902), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n562), .B(new_n387), .C1(new_n484), .C2(new_n485), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n659), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT34), .B(G104), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  NAND2_X1  g490(.A1(new_n552), .A2(new_n538), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n586), .A3(new_n591), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n561), .B(KEYINPUT102), .Z(new_n679));
  OAI211_X1 g493(.A(new_n387), .B(new_n679), .C1(new_n484), .C2(new_n485), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n659), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT104), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G9));
  NAND2_X1  g499(.A1(new_n242), .A2(new_n244), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(KEYINPUT36), .B2(new_n245), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n245), .A2(KEYINPUT36), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n242), .A2(new_n244), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n259), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n640), .B(new_n639), .C1(new_n646), .C2(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n656), .A2(new_n691), .A3(new_n486), .ZN(new_n692));
  INV_X1    g506(.A(new_n592), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  NOR2_X1   g510(.A1(new_n691), .A2(new_n486), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n385), .B1(new_n650), .B2(KEYINPUT32), .ZN(new_n698));
  INV_X1    g512(.A(G900), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n559), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n556), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n678), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n697), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  INV_X1    g519(.A(new_n641), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n701), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n709));
  INV_X1    g523(.A(new_n690), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n255), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n663), .A2(new_n586), .ZN(new_n712));
  INV_X1    g526(.A(new_n387), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT38), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n484), .B2(new_n485), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n453), .A2(new_n480), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n482), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n453), .A2(new_n480), .A3(new_n483), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(KEYINPUT38), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n708), .A2(KEYINPUT40), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n709), .A2(new_n714), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n382), .A2(new_n268), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n247), .B1(new_n373), .B2(new_n267), .ZN(new_n725));
  OAI21_X1  g539(.A(G472), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n365), .A2(new_n370), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n727), .B(new_n728), .C1(new_n650), .C2(KEYINPUT32), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT106), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n281), .ZN(G45));
  XOR2_X1   g546(.A(new_n667), .B(KEYINPUT33), .Z(new_n733));
  AOI22_X1  g547(.A1(new_n733), .A2(new_n669), .B1(new_n581), .B2(new_n665), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n702), .B(new_n734), .C1(new_n553), .C2(new_n591), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n697), .A2(new_n698), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  NOR2_X1   g551(.A1(new_n673), .A2(new_n672), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n646), .A2(new_n260), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n630), .A2(new_n631), .ZN(new_n740));
  OAI21_X1  g554(.A(G469), .B1(new_n740), .B2(G902), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n640), .A3(new_n632), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n738), .A2(new_n698), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NOR2_X1   g560(.A1(new_n680), .A2(new_n678), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(new_n698), .A3(new_n739), .A4(new_n743), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NOR2_X1   g563(.A1(new_n486), .A2(new_n742), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n698), .A2(new_n750), .A3(new_n693), .A4(new_n711), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NAND3_X1  g566(.A1(new_n255), .A2(KEYINPUT107), .A3(new_n261), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n646), .B2(new_n260), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n267), .B1(new_n374), .B2(new_n340), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n366), .B(new_n247), .C1(new_n363), .C2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n655), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n663), .A2(new_n586), .A3(new_n679), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n756), .A2(new_n750), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NAND2_X1  g577(.A1(new_n655), .A2(new_n758), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n646), .A2(new_n690), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n735), .A3(new_n750), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  NAND2_X1  g582(.A1(new_n756), .A2(new_n698), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n636), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n610), .A2(new_n614), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .A3(G469), .A4(new_n633), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n637), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n609), .A2(new_n615), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT83), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n609), .A2(new_n623), .A3(new_n615), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n601), .ZN(new_n778));
  INV_X1    g592(.A(new_n631), .ZN(new_n779));
  AOI211_X1 g593(.A(G469), .B(G902), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT109), .B(new_n640), .C1(new_n774), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n484), .A2(new_n485), .A3(new_n713), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n640), .B1(new_n774), .B2(new_n780), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n735), .A2(new_n781), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT42), .B1(new_n769), .B2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n782), .A2(new_n785), .A3(new_n781), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n663), .A2(new_n671), .A3(new_n701), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(KEYINPUT42), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n386), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n310), .ZN(G33));
  NAND3_X1  g607(.A1(new_n788), .A2(new_n386), .A3(new_n703), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n651), .B2(new_n765), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n656), .A2(KEYINPUT110), .A3(new_n711), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n663), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n671), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n663), .A2(KEYINPUT43), .A3(new_n734), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n782), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n802), .A2(new_n803), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n797), .B2(new_n798), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT112), .B1(new_n810), .B2(KEYINPUT44), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n805), .A2(new_n812), .A3(new_n806), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n807), .A2(KEYINPUT111), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n620), .A2(KEYINPUT45), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n620), .A2(KEYINPUT45), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(G469), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n637), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n780), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(KEYINPUT46), .A3(new_n637), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n823), .A2(new_n640), .A3(new_n707), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n808), .A2(new_n814), .A3(new_n815), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G137), .ZN(G39));
  AOI21_X1  g640(.A(KEYINPUT47), .B1(new_n823), .B2(new_n640), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  INV_X1    g642(.A(new_n640), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n828), .B(new_n829), .C1(new_n821), .C2(new_n822), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n370), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n375), .A2(new_n247), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n339), .A2(new_n342), .ZN(new_n834));
  INV_X1    g648(.A(new_n332), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n267), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n358), .A2(new_n338), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT29), .B1(new_n837), .B2(new_n268), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n833), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n649), .A2(new_n832), .B1(new_n839), .B2(new_n366), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n368), .B2(new_n367), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n262), .A3(new_n735), .A4(new_n782), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n831), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n201), .ZN(G42));
  INV_X1    g658(.A(new_n730), .ZN(new_n845));
  INV_X1    g659(.A(new_n801), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n756), .A3(new_n387), .A4(new_n640), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n741), .A2(new_n632), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(KEYINPUT113), .B1(KEYINPUT49), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT113), .B2(new_n847), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT114), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(KEYINPUT49), .ZN(new_n852));
  OR4_X1    g666(.A1(new_n845), .A2(new_n851), .A3(new_n721), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n764), .B1(new_n755), .B2(new_n753), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n804), .A2(new_n557), .A3(new_n750), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n782), .A2(new_n743), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT120), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n857), .A2(new_n557), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n739), .A3(new_n730), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n554), .B(new_n855), .C1(new_n860), .C2(new_n672), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n804), .A2(new_n557), .A3(new_n857), .A4(new_n858), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT48), .B1(new_n863), .B2(new_n769), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT48), .ZN(new_n865));
  INV_X1    g679(.A(new_n769), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n859), .A2(new_n865), .A3(new_n866), .A4(new_n804), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(KEYINPUT122), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n870));
  INV_X1    g684(.A(new_n868), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n861), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n721), .A2(new_n387), .A3(new_n742), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n804), .A2(new_n873), .A3(new_n557), .A4(new_n854), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT50), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n845), .A2(new_n262), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n800), .A3(new_n859), .A4(new_n734), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n859), .A2(new_n766), .A3(new_n804), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n741), .A2(new_n829), .A3(new_n632), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n831), .A2(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n557), .A2(new_n804), .A3(new_n854), .A4(new_n782), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n876), .A2(new_n878), .A3(new_n879), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n869), .A2(new_n872), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n876), .A2(new_n878), .A3(new_n889), .A4(new_n879), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n831), .A2(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n881), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n831), .A2(KEYINPUT119), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n883), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n888), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n886), .B1(new_n895), .B2(new_n880), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n744), .A2(new_n762), .A3(new_n751), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n591), .B(new_n587), .C1(new_n660), .C2(new_n662), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n671), .B1(new_n553), .B2(new_n591), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n680), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n653), .A2(new_n657), .A3(new_n902), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n692), .A2(new_n693), .B1(new_n386), .B2(new_n642), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n898), .A2(new_n748), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n759), .A2(new_n711), .A3(new_n735), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n782), .A2(new_n785), .A3(new_n781), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n584), .A2(new_n585), .A3(new_n701), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n589), .B2(new_n590), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n677), .A2(new_n909), .A3(KEYINPUT115), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT115), .B1(new_n677), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n706), .A3(new_n782), .A4(new_n711), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n906), .A2(new_n907), .B1(new_n913), .B2(new_n841), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n915), .A2(new_n787), .A3(new_n791), .A4(new_n794), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n897), .B1(new_n905), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n904), .A2(new_n903), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n744), .A2(new_n748), .A3(new_n762), .A4(new_n751), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n764), .A2(new_n789), .A3(new_n765), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n788), .ZN(new_n922));
  INV_X1    g736(.A(new_n691), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n698), .A2(new_n923), .A3(new_n782), .A4(new_n912), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n794), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n792), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n920), .A2(new_n926), .A3(KEYINPUT116), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n712), .A2(new_n486), .ZN(new_n928));
  NOR4_X1   g742(.A1(new_n783), .A2(new_n646), .A3(new_n690), .A4(new_n702), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n729), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n704), .A2(new_n767), .A3(new_n736), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT52), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n917), .A2(new_n927), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT53), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n903), .A2(new_n643), .A3(new_n694), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n744), .A2(new_n748), .A3(new_n762), .A4(new_n751), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n788), .A2(new_n698), .A3(new_n735), .A4(new_n756), .ZN(new_n940));
  AOI21_X1  g754(.A(G902), .B1(new_n349), .B2(new_n364), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT32), .B1(new_n941), .B2(new_n366), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n739), .B1(new_n942), .B2(new_n840), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n907), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n940), .A2(KEYINPUT42), .B1(new_n944), .B2(new_n790), .ZN(new_n945));
  INV_X1    g759(.A(new_n703), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n943), .A2(new_n907), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n914), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n938), .A2(new_n939), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  AOI22_X1  g763(.A1(new_n949), .A2(new_n897), .B1(new_n934), .B2(new_n933), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n927), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n937), .A2(KEYINPUT54), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n936), .A2(new_n951), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT54), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n711), .A3(new_n743), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n841), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n760), .A2(new_n486), .A3(new_n742), .ZN(new_n959));
  AOI22_X1  g773(.A1(new_n958), .A2(new_n693), .B1(new_n854), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT118), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n744), .A4(new_n748), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n904), .A2(KEYINPUT53), .A3(new_n903), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n919), .A2(KEYINPUT118), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n926), .A2(new_n962), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n931), .B(KEYINPUT52), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n954), .A2(new_n955), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n896), .A2(new_n953), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(G952), .A2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n853), .B1(new_n970), .B2(new_n971), .ZN(G75));
  NOR2_X1   g786(.A1(new_n216), .A2(G952), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n967), .B1(new_n936), .B2(new_n951), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(new_n247), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT56), .B1(new_n976), .B2(new_n482), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n442), .A2(new_n448), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n446), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT55), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n974), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  AOI211_X1 g796(.A(KEYINPUT56), .B(new_n980), .C1(new_n976), .C2(new_n482), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(G51));
  INV_X1    g798(.A(new_n740), .ZN(new_n985));
  INV_X1    g799(.A(new_n951), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n950), .B2(new_n927), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT54), .B1(new_n987), .B2(new_n967), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n969), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n637), .B(KEYINPUT57), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OR3_X1    g805(.A1(new_n975), .A2(new_n247), .A3(new_n818), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n973), .B1(new_n991), .B2(new_n992), .ZN(G54));
  NAND3_X1  g807(.A1(new_n976), .A2(KEYINPUT58), .A3(G475), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n973), .B1(new_n994), .B2(new_n550), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n976), .A2(KEYINPUT58), .A3(G475), .A4(new_n547), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(G60));
  NAND2_X1  g811(.A1(G478), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT59), .Z(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(new_n953), .B2(new_n969), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n974), .B1(new_n1000), .B2(new_n733), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n988), .A2(new_n969), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n668), .A2(new_n999), .ZN(new_n1003));
  AOI21_X1  g817(.A(KEYINPUT123), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1003), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n1005), .B(new_n1006), .C1(new_n988), .C2(new_n969), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1001), .A2(new_n1004), .A3(new_n1007), .ZN(G63));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT60), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n256), .B1(new_n975), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n687), .A2(new_n689), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1010), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1012), .B(new_n1013), .C1(new_n987), .C2(new_n967), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1011), .A2(new_n974), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT124), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT61), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1013), .B1(new_n987), .B2(new_n967), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n973), .B1(new_n1021), .B2(new_n256), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1022), .A2(new_n1017), .A3(new_n1018), .A4(new_n1014), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1020), .A2(new_n1023), .ZN(G66));
  INV_X1    g838(.A(G224), .ZN(new_n1025));
  OAI21_X1  g839(.A(G953), .B1(new_n560), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n920), .B2(G953), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n978), .B1(G898), .B2(new_n216), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G69));
  XNOR2_X1  g843(.A(new_n381), .B(new_n531), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n704), .A2(new_n767), .A3(new_n736), .ZN(new_n1031));
  OR3_X1    g845(.A1(new_n731), .A2(KEYINPUT62), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n782), .A2(new_n706), .A3(new_n707), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1033), .A2(new_n900), .A3(new_n901), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n843), .B1(new_n386), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(KEYINPUT62), .B1(new_n731), .B2(new_n1031), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(new_n825), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1030), .B1(new_n1038), .B2(new_n216), .ZN(new_n1039));
  INV_X1    g853(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(G953), .B1(new_n612), .B2(new_n699), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(KEYINPUT125), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n824), .A2(new_n866), .A3(new_n928), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1043), .B(new_n794), .C1(new_n831), .C2(new_n842), .ZN(new_n1044));
  NOR3_X1   g858(.A1(new_n1044), .A2(new_n792), .A3(new_n1031), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n825), .A2(new_n216), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1030), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1047), .B1(G900), .B2(G953), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OR2_X1    g863(.A1(new_n1041), .A2(KEYINPUT125), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1040), .A2(new_n1042), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1049), .ZN(new_n1052));
  OAI211_X1 g866(.A(KEYINPUT125), .B(new_n1041), .C1(new_n1052), .C2(new_n1039), .ZN(new_n1053));
  AND2_X1   g867(.A1(new_n1051), .A2(new_n1053), .ZN(G72));
  NAND2_X1  g868(.A1(G472), .A2(G902), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT63), .Z(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1038), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1057), .B1(new_n1058), .B2(new_n920), .ZN(new_n1059));
  INV_X1    g873(.A(new_n724), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n937), .A2(new_n952), .ZN(new_n1061));
  NOR2_X1   g875(.A1(new_n837), .A2(new_n267), .ZN(new_n1062));
  OR3_X1    g876(.A1(new_n724), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  OAI22_X1  g877(.A1(new_n1059), .A2(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n815), .A2(new_n814), .ZN(new_n1065));
  OAI21_X1  g879(.A(new_n824), .B1(new_n807), .B2(KEYINPUT111), .ZN(new_n1066));
  OAI211_X1 g880(.A(new_n1045), .B(new_n920), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT126), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1067), .A2(new_n1068), .A3(new_n1056), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1069), .A2(new_n1062), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1068), .B1(new_n1067), .B2(new_n1056), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n974), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g886(.A(KEYINPUT127), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g888(.A(KEYINPUT127), .B(new_n974), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(G57));
endmodule


