//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  AND2_X1   g000(.A1(G127gat), .A2(G134gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR3_X1   g004(.A1(new_n205), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G120gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n205), .A2(G113gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n207), .A2(new_n209), .B1(new_n204), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n216), .A2(KEYINPUT26), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n216), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT27), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G183gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n225), .A2(G183gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n223), .A2(KEYINPUT27), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT69), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT69), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(G190gat), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n229), .B1(new_n235), .B2(new_n227), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n224), .A2(new_n226), .A3(new_n233), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n224), .B2(new_n226), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n228), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT28), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT70), .A3(new_n229), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n222), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  INV_X1    g045(.A(G176gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT23), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n218), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n223), .A2(new_n228), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT65), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n254), .A4(new_n255), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n248), .A2(new_n245), .A3(new_n249), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n253), .A2(new_n258), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  INV_X1    g065(.A(new_n252), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT66), .B1(new_n216), .B2(KEYINPUT23), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(KEYINPUT25), .A3(new_n262), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n271), .A2(new_n272), .A3(new_n256), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  AND4_X1   g073(.A1(new_n218), .A2(new_n262), .A3(new_n268), .A4(new_n251), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n257), .A2(KEYINPUT67), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(new_n254), .A3(new_n255), .A4(new_n270), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n275), .A2(KEYINPUT68), .A3(KEYINPUT25), .A4(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n265), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n215), .B1(new_n244), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n222), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT70), .B1(new_n242), .B2(new_n229), .ZN(new_n282));
  INV_X1    g081(.A(new_n229), .ZN(new_n283));
  AOI211_X1 g082(.A(new_n237), .B(new_n283), .C1(new_n241), .C2(KEYINPUT28), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n207), .A2(new_n209), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n214), .A2(new_n204), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n274), .A3(new_n278), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT64), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n280), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(G71gat), .B(G99gat), .Z(new_n294));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT33), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n293), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n297), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n303));
  INV_X1    g102(.A(new_n293), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n303), .B(new_n296), .C1(new_n304), .C2(KEYINPUT33), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT34), .ZN(new_n307));
  INV_X1    g106(.A(new_n292), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(KEYINPUT73), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n280), .A2(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  AOI211_X1 g111(.A(new_n292), .B(new_n309), .C1(new_n280), .C2(new_n290), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n302), .A2(new_n305), .A3(new_n314), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n318));
  XOR2_X1   g117(.A(G197gat), .B(G204gat), .Z(new_n319));
  AOI21_X1  g118(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT79), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n322), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT74), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n318), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G155gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G162gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G148gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(G141gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n335), .A2(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n334), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT76), .B(G162gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT2), .B1(new_n343), .B2(new_n332), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346));
  INV_X1    g145(.A(G141gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G148gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n340), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n334), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n326), .A2(new_n323), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n342), .A2(new_n344), .B1(new_n349), .B2(new_n334), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n328), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n318), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n328), .B1(new_n353), .B2(KEYINPUT29), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n351), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n362), .A2(G228gat), .A3(G233gat), .A4(new_n357), .ZN(new_n363));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G22gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(KEYINPUT80), .A2(G22gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n366), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n360), .A2(new_n363), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n360), .B2(new_n363), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n316), .A2(new_n317), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n244), .B2(new_n279), .ZN(new_n382));
  INV_X1    g181(.A(new_n353), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n285), .B2(new_n289), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n381), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n318), .B1(new_n244), .B2(new_n279), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n380), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n388), .B2(new_n382), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n379), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n382), .B1(new_n384), .B2(new_n381), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n353), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n378), .A3(new_n385), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(KEYINPUT30), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n392), .A2(new_n395), .A3(new_n378), .A4(new_n385), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n354), .A2(new_n215), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n354), .A2(new_n215), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n215), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n355), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n351), .A2(new_n288), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n398), .ZN(new_n409));
  INV_X1    g208(.A(new_n405), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n400), .B1(new_n354), .B2(new_n215), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(KEYINPUT77), .B2(new_n401), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n404), .B(new_n413), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G1gat), .B(G29gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n418), .ZN(new_n428));
  INV_X1    g227(.A(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n423), .A2(KEYINPUT78), .A3(new_n424), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n397), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT35), .B1(new_n375), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n302), .A2(new_n305), .A3(new_n314), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n314), .B1(new_n302), .B2(new_n305), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n401), .A2(KEYINPUT77), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n399), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(new_n416), .B1(new_n355), .B2(new_n403), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n443), .A2(new_n413), .B1(new_n406), .B2(new_n411), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n422), .B(KEYINPUT81), .Z(new_n445));
  OAI211_X1 g244(.A(new_n423), .B(new_n424), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n440), .B1(new_n446), .B2(new_n433), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n439), .A2(new_n397), .A3(new_n374), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n436), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n437), .B2(new_n438), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n316), .A2(KEYINPUT36), .A3(new_n317), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n374), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n444), .A2(new_n445), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n408), .A2(new_n398), .A3(new_n405), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n458), .A2(KEYINPUT39), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n443), .B2(new_n405), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n404), .B1(new_n415), .B2(new_n417), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n410), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n445), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n456), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n457), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n394), .A2(new_n396), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n446), .A2(new_n393), .A3(new_n433), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT37), .B1(new_n386), .B2(new_n389), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n392), .A2(new_n471), .A3(new_n385), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n379), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n392), .A2(new_n385), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n378), .B1(new_n475), .B2(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n470), .B1(new_n476), .B2(new_n472), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n467), .B(new_n374), .C1(new_n474), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n455), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n449), .A2(new_n479), .A3(KEYINPUT84), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT84), .B1(new_n449), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT98), .ZN(new_n483));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G78gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(KEYINPUT21), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT94), .ZN(new_n490));
  XOR2_X1   g289(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G183gat), .B(G211gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G1gat), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT92), .C1(G1gat), .C2(new_n495), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT93), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(KEYINPUT21), .B2(new_n488), .ZN(new_n502));
  XNOR2_X1  g301(.A(G127gat), .B(G155gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(G231gat), .A2(G233gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n502), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n494), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G43gat), .B(G50gat), .Z(new_n508));
  INV_X1    g307(.A(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n510), .A2(KEYINPUT15), .A3(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT88), .B(G36gat), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G29gat), .ZN(new_n515));
  NOR3_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(KEYINPUT87), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n515), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(KEYINPUT89), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT89), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n516), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n510), .A2(KEYINPUT15), .A3(new_n512), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n515), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n523), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT91), .B1(new_n535), .B2(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n522), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n528), .B(KEYINPUT90), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(new_n533), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n536), .A2(new_n542), .B1(KEYINPUT17), .B2(new_n535), .ZN(new_n543));
  XOR2_X1   g342(.A(G99gat), .B(G106gat), .Z(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G99gat), .ZN(new_n546));
  INV_X1    g345(.A(G106gat), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT8), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(G85gat), .B2(G92gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT96), .ZN(new_n552));
  NOR2_X1   g351(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n549), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n551), .A2(KEYINPUT96), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(KEYINPUT96), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n545), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n545), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G190gat), .B(G218gat), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n562), .A2(new_n535), .ZN(new_n566));
  AND2_X1   g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(KEYINPUT41), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n565), .B1(new_n563), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n567), .A2(KEYINPUT41), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n569), .A2(new_n570), .B1(KEYINPUT97), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n563), .A2(new_n568), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n564), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n573), .B(KEYINPUT97), .Z(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n507), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n543), .A2(new_n500), .B1(new_n539), .B2(new_n501), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT18), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n536), .A2(new_n542), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n500), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n501), .A2(new_n539), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(KEYINPUT18), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n500), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n535), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n584), .B(KEYINPUT13), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT85), .B1(new_n585), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(G197gat), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT11), .B(G169gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT12), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT85), .B(new_n605), .C1(new_n597), .C2(new_n585), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n488), .ZN(new_n608));
  INV_X1    g407(.A(new_n561), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n559), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n560), .A2(new_n488), .A3(new_n561), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n560), .A2(KEYINPUT10), .A3(new_n488), .A4(new_n561), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G230gat), .ZN(new_n616));
  INV_X1    g415(.A(G233gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  AND2_X1   g422(.A1(new_n610), .A2(new_n611), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n620), .B(new_n623), .C1(new_n624), .C2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n619), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n618), .B1(new_n613), .B2(new_n614), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n582), .A2(new_n607), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n482), .A2(new_n483), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n449), .A2(new_n479), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT84), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n449), .A2(new_n479), .A3(KEYINPUT84), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n434), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT99), .B(G1gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1324gat));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644));
  INV_X1    g443(.A(new_n397), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n483), .B1(new_n482), .B2(new_n631), .ZN(new_n646));
  AND4_X1   g445(.A1(new_n483), .A2(new_n635), .A3(new_n636), .A4(new_n631), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(G8gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n639), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n644), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n397), .B(new_n650), .C1(new_n632), .C2(new_n638), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT100), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n499), .B1(new_n639), .B2(new_n645), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n657), .B2(new_n654), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n652), .A2(new_n644), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n656), .A2(new_n661), .ZN(G1325gat));
  INV_X1    g461(.A(new_n639), .ZN(new_n663));
  INV_X1    g462(.A(new_n439), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n663), .A2(G15gat), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n663), .B2(new_n453), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n639), .A2(new_n454), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(KEYINPUT101), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(G1327gat));
  NAND2_X1  g475(.A1(new_n449), .A2(KEYINPUT104), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n436), .A2(new_n678), .A3(new_n448), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n396), .A2(new_n394), .B1(new_n432), .B2(new_n433), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n682), .B2(new_n374), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n435), .A2(KEYINPUT102), .A3(new_n454), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n453), .A2(new_n478), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n685), .A2(KEYINPUT103), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n453), .A2(new_n478), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n684), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n680), .B1(new_n687), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n575), .A2(new_n580), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n694));
  NAND3_X1  g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n635), .A2(new_n636), .A3(new_n693), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n607), .A2(new_n507), .A3(new_n630), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n434), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n482), .A2(new_n693), .A3(new_n699), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n702), .A2(G29gat), .A3(new_n434), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(KEYINPUT45), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(G1328gat));
  OAI21_X1  g505(.A(new_n514), .B1(new_n700), .B2(new_n397), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n397), .A2(new_n514), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT46), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  OR3_X1    g508(.A1(new_n702), .A2(KEYINPUT46), .A3(new_n708), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  NOR2_X1   g510(.A1(new_n664), .A2(G43gat), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n702), .A2(new_n713), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n714));
  INV_X1    g513(.A(new_n453), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n715), .A3(new_n699), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1330gat));
  NOR3_X1   g518(.A1(new_n702), .A2(G50gat), .A3(new_n374), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n454), .A3(new_n699), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(G50gat), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT48), .ZN(G1331gat));
  OAI21_X1  g522(.A(KEYINPUT103), .B1(new_n685), .B2(new_n686), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n689), .A2(new_n688), .A3(new_n690), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n724), .A2(new_n725), .B1(new_n677), .B2(new_n679), .ZN(new_n726));
  INV_X1    g525(.A(new_n607), .ZN(new_n727));
  INV_X1    g526(.A(new_n630), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n582), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n640), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT107), .B(G57gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1332gat));
  AOI21_X1  g534(.A(new_n397), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT109), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n732), .A2(new_n715), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n664), .A2(G71gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(G71gat), .B1(new_n732), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n732), .A2(new_n454), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(G78gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  INV_X1    g547(.A(new_n507), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n729), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n698), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n434), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n727), .A2(new_n507), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n692), .A2(new_n693), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT51), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n692), .A2(new_n757), .A3(new_n693), .A4(new_n754), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n630), .A3(new_n758), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n434), .A2(G85gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n753), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(new_n694), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n726), .A2(new_n581), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n482), .B2(new_n693), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n645), .B(new_n751), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n750), .B1(new_n695), .B2(new_n697), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(KEYINPUT111), .A3(new_n645), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(G92gat), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n397), .A2(G92gat), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n756), .A2(new_n630), .A3(new_n758), .A4(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(G92gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n769), .B2(new_n645), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n752), .B2(new_n453), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n439), .A2(new_n546), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n759), .B2(new_n783), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n752), .B2(new_n374), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n374), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(new_n786), .C1(new_n759), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n759), .A2(new_n788), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n547), .B1(new_n769), .B2(new_n454), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1339gat));
  NAND3_X1  g592(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n620), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n623), .B1(new_n628), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  INV_X1    g598(.A(new_n625), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n604), .A2(new_n801), .A3(new_n606), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT112), .B1(new_n594), .B2(new_n595), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n804));
  INV_X1    g603(.A(new_n595), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n589), .A2(new_n593), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n583), .A2(new_n584), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n602), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n588), .A2(new_n584), .A3(new_n589), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT18), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(new_n590), .A3(new_n596), .A4(new_n605), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n813), .A3(new_n630), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n693), .B1(new_n802), .B2(new_n814), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n693), .A2(new_n801), .A3(new_n813), .A4(new_n809), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n749), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n730), .A2(new_n607), .A3(new_n728), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n640), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n645), .A3(new_n375), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n727), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n211), .A2(KEYINPUT113), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n211), .A2(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n630), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n507), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G127gat), .ZN(G1342gat));
  INV_X1    g629(.A(new_n821), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n831), .B2(new_n581), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n693), .A2(new_n397), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT114), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n375), .A2(G134gat), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n640), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n809), .A2(new_n813), .A3(new_n840), .A4(new_n630), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n814), .A2(KEYINPUT115), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n802), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n816), .B1(new_n843), .B2(new_n581), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n818), .B1(new_n844), .B2(new_n507), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n454), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n453), .A2(new_n640), .A3(new_n397), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n374), .B1(new_n817), .B2(new_n818), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n727), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n839), .B1(new_n852), .B2(G141gat), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n819), .A2(new_n640), .A3(new_n454), .A4(new_n453), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n727), .A2(new_n347), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n645), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n852), .B2(G141gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n853), .A2(new_n857), .A3(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  AOI221_X4 g658(.A(new_n856), .B1(new_n839), .B2(new_n859), .C1(new_n852), .C2(G141gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n858), .A2(new_n860), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n854), .A2(new_n645), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n336), .A2(new_n338), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n630), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n849), .A2(KEYINPUT57), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n845), .B2(new_n454), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n848), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n630), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n865), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n847), .A2(new_n851), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT59), .B(new_n863), .C1(new_n872), .C2(new_n630), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n864), .B1(new_n871), .B2(new_n873), .ZN(G1345gat));
  NOR3_X1   g673(.A1(new_n854), .A2(new_n645), .A3(new_n749), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g675(.A(G155gat), .B1(new_n875), .B2(KEYINPUT117), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n749), .A2(new_n332), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n876), .A2(new_n877), .B1(new_n872), .B2(new_n878), .ZN(G1346gat));
  AND2_X1   g678(.A1(new_n872), .A2(new_n693), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n834), .A2(new_n343), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n880), .A2(new_n343), .B1(new_n854), .B2(new_n881), .ZN(G1347gat));
  NAND2_X1  g681(.A1(new_n645), .A2(new_n434), .ZN(new_n883));
  OR3_X1    g682(.A1(new_n664), .A2(new_n883), .A3(KEYINPUT118), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT118), .B1(new_n664), .B2(new_n883), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n454), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n819), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n246), .A3(new_n607), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n640), .B1(new_n817), .B2(new_n818), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n375), .A2(new_n397), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n727), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n888), .B1(new_n893), .B2(new_n246), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n887), .B2(new_n728), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n630), .A2(new_n247), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n891), .B2(new_n896), .ZN(G1349gat));
  NOR2_X1   g696(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n898));
  AND2_X1   g697(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n749), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT119), .B1(new_n887), .B2(new_n749), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(G183gat), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n892), .B(new_n507), .C1(new_n239), .C2(new_n240), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n898), .B(new_n899), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  AND4_X1   g703(.A1(KEYINPUT120), .A2(new_n902), .A3(KEYINPUT60), .A4(new_n903), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1350gat));
  NOR3_X1   g705(.A1(new_n891), .A2(G190gat), .A3(new_n581), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT121), .ZN(new_n908));
  OAI21_X1  g707(.A(G190gat), .B1(new_n887), .B2(new_n581), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(KEYINPUT122), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n908), .A2(new_n912), .A3(new_n914), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n715), .A2(new_n397), .A3(new_n374), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n889), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n727), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n715), .A2(new_n883), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT123), .Z(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n868), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n727), .A2(G197gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  NAND3_X1  g724(.A1(new_n868), .A2(new_n922), .A3(new_n630), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G204gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n917), .A2(G204gat), .A3(new_n728), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT62), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1353gat));
  AND2_X1   g729(.A1(new_n921), .A2(new_n507), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n866), .A2(new_n867), .ZN(new_n933));
  OAI21_X1  g732(.A(G211gat), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT63), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(KEYINPUT63), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n917), .A2(G211gat), .A3(new_n749), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT125), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(G1354gat));
  AOI21_X1  g738(.A(G218gat), .B1(new_n918), .B2(new_n693), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n693), .A2(G218gat), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT126), .Z(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n923), .B2(new_n942), .ZN(G1355gat));
endmodule


