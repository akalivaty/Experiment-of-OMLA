//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n202), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT64), .B(G238), .Z(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n223), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n226), .B(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n221), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT66), .B(G250), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT14), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G226), .A2(G1698), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(new_n207), .B2(G1698), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(KEYINPUT71), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT71), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n252), .A2(new_n253), .B1(G33), .B2(G97), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n259), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n259), .A2(new_n266), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G238), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n261), .A2(new_n264), .A3(new_n269), .A4(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n250), .B1(new_n276), .B2(G169), .ZN(new_n277));
  INV_X1    g0077(.A(G169), .ZN(new_n278));
  AOI211_X1 g0078(.A(KEYINPUT14), .B(new_n278), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  INV_X1    g0083(.A(G20), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n283), .A2(new_n284), .A3(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n223), .B2(new_n257), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT67), .B1(new_n265), .B2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n290), .A2(new_n284), .A3(G1), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n288), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G68), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n284), .A2(new_n257), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n284), .A2(G33), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n294), .A2(new_n202), .B1(new_n295), .B2(new_n213), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n284), .A2(G68), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT11), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n283), .A2(G1), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n297), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT12), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n293), .A2(new_n300), .A3(new_n301), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n282), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n276), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n274), .B2(new_n275), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n203), .A2(G20), .ZN(new_n314));
  INV_X1    g0114(.A(G150), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n315), .B2(new_n294), .C1(new_n316), .C2(new_n295), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n287), .B1(new_n202), .B2(new_n285), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n292), .A2(G50), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G223), .A2(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G222), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n253), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(new_n260), .C1(G77), .C2(new_n253), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n271), .A2(G226), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n269), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n320), .A2(new_n321), .B1(new_n328), .B2(new_n308), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT9), .B1(new_n318), .B2(new_n319), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT10), .ZN(new_n334));
  INV_X1    g0134(.A(new_n328), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n320), .B1(new_n335), .B2(G169), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(G179), .C2(new_n328), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G20), .A2(G77), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT15), .B(G87), .Z(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(new_n316), .B(KEYINPUT69), .Z(new_n345));
  OAI221_X1 g0145(.A(new_n342), .B1(new_n295), .B2(new_n344), .C1(new_n345), .C2(new_n294), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n287), .B1(new_n213), .B2(new_n285), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n292), .A2(G77), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n323), .A2(G232), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n253), .B(new_n349), .C1(new_n219), .C2(new_n323), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n260), .C1(G107), .C2(new_n253), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n268), .B1(new_n271), .B2(G244), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G190), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n352), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n347), .A2(new_n348), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n313), .A2(new_n341), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT7), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT72), .B(G33), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n363), .B2(G20), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n358), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT73), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G33), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n360), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(new_n365), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n364), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G68), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n294), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n206), .A2(new_n218), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n379), .A2(new_n201), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n380), .B2(G20), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n360), .A2(new_n383), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n284), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n384), .A2(new_n365), .B1(new_n386), .B2(new_n358), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n381), .B1(new_n387), .B2(new_n218), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n287), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n212), .A2(G1698), .ZN(new_n394));
  OR2_X1    g0194(.A1(G223), .A2(G1698), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n371), .A2(new_n394), .A3(new_n360), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n268), .B1(new_n398), .B2(new_n260), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n270), .A2(new_n207), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT75), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n259), .B1(new_n396), .B2(new_n397), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT75), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n400), .A4(new_n268), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n310), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n398), .A2(new_n260), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n401), .A3(new_n269), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n406), .B1(G190), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n287), .ZN(new_n410));
  INV_X1    g0210(.A(new_n381), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n375), .B2(G68), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT74), .A3(new_n390), .ZN(new_n414));
  INV_X1    g0214(.A(new_n316), .ZN(new_n415));
  MUX2_X1   g0215(.A(new_n285), .B(new_n292), .S(new_n415), .Z(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n393), .A2(new_n409), .A3(new_n414), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n278), .B1(new_n402), .B2(new_n405), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n408), .A2(G179), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n423), .B2(new_n426), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n393), .A2(new_n417), .A3(new_n414), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n429), .A2(KEYINPUT18), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT18), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n420), .B(new_n422), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n354), .A2(G179), .ZN(new_n435));
  XOR2_X1   g0235(.A(new_n435), .B(KEYINPUT70), .Z(new_n436));
  NAND2_X1  g0236(.A1(new_n354), .A2(new_n278), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n347), .A2(new_n348), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n357), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G20), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n287), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n284), .C1(G33), .C2(new_n220), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT20), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n287), .A3(new_n443), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT20), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT80), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n450), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n302), .A2(G20), .A3(new_n442), .ZN(new_n454));
  AOI211_X1 g0254(.A(new_n287), .B(new_n285), .C1(new_n265), .C2(G33), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G116), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n323), .A2(G264), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n221), .A2(new_n323), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n371), .A2(new_n360), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n385), .A2(G303), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n259), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n265), .A2(G45), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT77), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT77), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n265), .A4(G45), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n471), .A2(G274), .A3(new_n259), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n466), .A2(new_n472), .A3(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G270), .A3(new_n259), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n463), .A2(new_n473), .A3(G190), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n457), .A2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n474), .A2(new_n267), .A3(new_n260), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n310), .B1(new_n479), .B2(new_n475), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n371), .A2(new_n284), .A3(G68), .A4(new_n360), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n284), .B1(new_n255), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n208), .A2(new_n220), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n484), .B1(new_n295), .B2(new_n220), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n491), .B(new_n484), .C1(new_n295), .C2(new_n220), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n483), .A2(new_n488), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n287), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n344), .A2(new_n285), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n455), .A2(new_n343), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(G238), .A2(G1698), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n214), .B2(G1698), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n371), .A3(new_n360), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n368), .A2(new_n370), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G116), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n259), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n465), .A2(new_n209), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n265), .A2(new_n267), .A3(G45), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n259), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n280), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n278), .B1(new_n503), .B2(new_n507), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n497), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n500), .A2(new_n502), .ZN(new_n512));
  OAI211_X1 g0312(.A(G190), .B(new_n506), .C1(new_n512), .C2(new_n259), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n493), .A2(new_n287), .B1(new_n285), .B2(new_n344), .ZN(new_n514));
  OAI21_X1  g0314(.A(G200), .B1(new_n503), .B2(new_n507), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n455), .A2(G87), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT79), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n511), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n482), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n285), .A2(new_n220), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n455), .A2(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n384), .A2(new_n365), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n386), .A2(new_n358), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n486), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n294), .A2(new_n213), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n220), .A2(new_n486), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n284), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n523), .B(new_n524), .C1(new_n535), .C2(new_n410), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n323), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n253), .B2(G250), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n446), .B(new_n537), .C1(new_n539), .C2(new_n323), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT4), .B1(new_n363), .B2(G244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n260), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n474), .A2(new_n259), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G257), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n544), .A3(new_n473), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n278), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n542), .A2(new_n544), .A3(new_n280), .A4(new_n473), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n536), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n528), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n532), .A2(new_n533), .ZN(new_n550));
  OAI221_X1 g0350(.A(new_n549), .B1(new_n550), .B2(new_n284), .C1(new_n387), .C2(new_n486), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n287), .B1(new_n220), .B2(new_n285), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n542), .A2(new_n544), .A3(G190), .A4(new_n473), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n524), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n501), .A2(new_n284), .A3(G116), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT23), .B1(new_n284), .B2(G107), .ZN(new_n559));
  OR3_X1    g0359(.A1(new_n284), .A2(KEYINPUT23), .A3(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n371), .A2(new_n284), .A3(G87), .A4(new_n360), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT81), .ZN(new_n566));
  OR4_X1    g0366(.A1(KEYINPUT22), .A2(new_n385), .A3(G20), .A4(new_n208), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n568), .A3(KEYINPUT22), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n563), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n287), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n455), .A2(G107), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n302), .A2(G20), .A3(new_n486), .ZN(new_n576));
  XOR2_X1   g0376(.A(new_n576), .B(KEYINPUT25), .Z(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n221), .A2(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n209), .A2(new_n323), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n371), .A2(new_n360), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n501), .A2(G294), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n259), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n543), .B2(G264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n473), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n278), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n280), .A3(new_n473), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n479), .A2(new_n475), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(G169), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT21), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n463), .A2(new_n473), .A3(G179), .A4(new_n475), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n457), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n585), .A2(new_n310), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G190), .B2(new_n585), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n574), .A2(new_n599), .A3(new_n575), .A4(new_n577), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n557), .A2(new_n588), .A3(new_n597), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n441), .A2(new_n601), .ZN(G372));
  INV_X1    g0402(.A(new_n339), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n312), .A2(new_n439), .ZN(new_n605));
  OR3_X1    g0405(.A1(new_n307), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n418), .B(KEYINPUT17), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n307), .B2(new_n605), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n429), .A2(new_n430), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n603), .B1(new_n615), .B2(new_n334), .ZN(new_n616));
  INV_X1    g0416(.A(new_n600), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n506), .B(KEYINPUT83), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n503), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n497), .B(new_n509), .C1(G169), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(G200), .B1(new_n618), .B2(new_n503), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n514), .A3(new_n513), .A4(new_n516), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n548), .A3(new_n555), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT84), .B1(new_n617), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n588), .A2(new_n597), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n548), .A2(new_n555), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT84), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n600), .A3(new_n630), .A4(new_n625), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n548), .A2(KEYINPUT26), .A3(new_n624), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n536), .A2(new_n546), .A3(new_n547), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n521), .A3(new_n519), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n621), .B(new_n633), .C1(KEYINPUT26), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n440), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n616), .A2(new_n638), .ZN(G369));
  NOR2_X1   g0439(.A1(new_n283), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n265), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n578), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n588), .B1(new_n647), .B2(new_n617), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n588), .A2(new_n646), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n597), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n649), .ZN(new_n656));
  INV_X1    g0456(.A(new_n653), .ZN(new_n657));
  INV_X1    g0457(.A(new_n646), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n457), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n597), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n481), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n656), .A2(new_n663), .ZN(G399));
  NOR2_X1   g0464(.A1(new_n487), .A2(G116), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT87), .Z(new_n666));
  INV_X1    g0466(.A(new_n227), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(G1), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT88), .Z(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n231), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT28), .ZN(new_n673));
  INV_X1    g0473(.A(new_n508), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n595), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n545), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT30), .A4(new_n584), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n584), .A2(new_n473), .A3(new_n544), .A4(new_n542), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n479), .A2(G179), .A3(new_n508), .A4(new_n475), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(G179), .B1(new_n479), .B2(new_n475), .ZN(new_n682));
  INV_X1    g0482(.A(new_n619), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n585), .A3(new_n545), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT31), .B1(new_n685), .B2(new_n646), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT89), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n646), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n685), .A2(KEYINPUT31), .A3(new_n646), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n511), .A2(new_n520), .A3(new_n517), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n520), .B1(new_n511), .B2(new_n517), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n697), .A3(new_n481), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n629), .A3(new_n600), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n628), .A2(new_n699), .A3(new_n646), .ZN(new_n700));
  OAI21_X1  g0500(.A(G330), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT90), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n688), .B(new_n694), .C1(new_n601), .C2(new_n646), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n556), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n548), .A2(new_n555), .A3(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n628), .A2(new_n711), .A3(new_n600), .A4(new_n623), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n620), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n634), .B2(new_n623), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n646), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT92), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n646), .B1(new_n632), .B2(new_n636), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n722), .A3(KEYINPUT29), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n707), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n673), .B1(new_n725), .B2(G1), .ZN(G364));
  AOI21_X1  g0526(.A(new_n265), .B1(new_n640), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n668), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n662), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n661), .A2(G330), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n253), .A2(G355), .A3(new_n227), .ZN(new_n734));
  INV_X1    g0534(.A(G45), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n245), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n363), .A2(new_n667), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G45), .B2(new_n231), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n734), .B1(G116), .B2(new_n227), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n286), .B1(G20), .B2(new_n278), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n743), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n284), .A2(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n377), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n284), .B1(new_n748), .B2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G97), .ZN(new_n754));
  NAND3_X1  g0554(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT94), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(G190), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n751), .B(new_n754), .C1(new_n202), .C2(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n757), .A2(new_n308), .A3(new_n758), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n760), .B1(G68), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n284), .A2(new_n308), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n310), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n280), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n747), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n763), .A2(new_n768), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(G77), .B1(new_n771), .B2(G58), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT93), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n764), .A2(new_n747), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n486), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n762), .A2(new_n253), .A3(new_n767), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n385), .B1(new_n752), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n749), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G322), .A2(new_n771), .B1(new_n781), .B2(G329), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n769), .ZN(new_n784));
  INV_X1    g0584(.A(new_n775), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n780), .B(new_n784), .C1(G283), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n759), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G326), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n766), .A2(G303), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT33), .B(G317), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n761), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n778), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n742), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n745), .B1(new_n746), .B2(new_n793), .C1(new_n661), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n733), .B1(new_n796), .B2(new_n730), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT96), .Z(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  NAND2_X1  g0599(.A1(new_n438), .A2(new_n646), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n356), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n439), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n439), .B2(new_n646), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n720), .A2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n646), .B(new_n803), .C1(new_n632), .C2(new_n636), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n707), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n707), .A2(KEYINPUT99), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n706), .A2(new_n805), .A3(new_n807), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n811), .A2(new_n730), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n761), .A2(G150), .B1(G143), .B2(new_n771), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n816), .B2(new_n759), .C1(new_n377), .C2(new_n769), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n363), .B1(new_n202), .B2(new_n765), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n775), .A2(new_n218), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G58), .C2(new_n753), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n818), .B(new_n821), .C1(new_n822), .C2(new_n749), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n775), .A2(new_n208), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(G311), .B2(new_n781), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(new_n771), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT97), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n385), .B1(new_n765), .B2(new_n486), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n754), .B1(new_n827), .B2(new_n779), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n761), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  INV_X1    g0632(.A(G303), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n759), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n830), .B(new_n834), .C1(new_n828), .C2(new_n829), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n826), .B(new_n835), .C1(new_n442), .C2(new_n769), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n746), .B1(new_n823), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n743), .A2(new_n740), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n213), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n839), .B(new_n729), .C1(new_n804), .C2(new_n741), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n814), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n412), .A2(KEYINPUT16), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n416), .B1(new_n843), .B2(new_n413), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n644), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n614), .B2(new_n607), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n408), .A2(new_n404), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n403), .A2(new_n400), .A3(new_n268), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT75), .ZN(new_n850));
  AOI21_X1  g0650(.A(G169), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT76), .B1(new_n851), .B2(new_n425), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n844), .B1(new_n854), .B2(new_n644), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n855), .B2(new_n421), .ZN(new_n856));
  INV_X1    g0656(.A(new_n644), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n430), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n610), .A2(new_n858), .A3(new_n859), .A4(new_n418), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n842), .B1(new_n847), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n433), .A2(new_n845), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT101), .B1(new_n691), .B2(KEYINPUT31), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n686), .B2(new_n687), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(new_n601), .C2(new_n646), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n305), .A2(new_n646), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n871), .B1(new_n311), .B2(new_n309), .C1(new_n282), .C2(new_n306), .ZN(new_n872));
  OR3_X1    g0672(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n305), .B(new_n646), .C1(new_n873), .C2(new_n312), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n870), .A2(new_n875), .A3(new_n804), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI221_X4 g0679(.A(new_n842), .B1(new_n856), .B2(new_n860), .C1(new_n433), .C2(new_n845), .ZN(new_n880));
  INV_X1    g0680(.A(new_n858), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n431), .A2(new_n432), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n422), .A2(new_n420), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n610), .A2(new_n858), .A3(new_n418), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n860), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT40), .B(new_n876), .C1(new_n880), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n440), .A2(new_n870), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n890), .B(new_n891), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(G330), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n439), .A2(new_n646), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n806), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n866), .A2(new_n875), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n880), .B2(new_n888), .ZN(new_n899));
  INV_X1    g0699(.A(new_n307), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n646), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n882), .A2(new_n644), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n440), .A2(new_n719), .A3(new_n721), .A4(new_n723), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n906), .A2(new_n616), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n893), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n265), .B2(new_n640), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT35), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n230), .B1(new_n550), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(G116), .C1(new_n911), .C2(new_n550), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n379), .A2(new_n231), .A3(new_n213), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT100), .Z(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(G50), .B2(new_n218), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n283), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n910), .A2(new_n914), .A3(new_n918), .ZN(G367));
  NAND2_X1  g0719(.A1(new_n536), .A2(new_n646), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n711), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n634), .A2(new_n646), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n653), .A2(new_n654), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT42), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n548), .B1(new_n921), .B2(new_n588), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n926), .A2(new_n927), .B1(new_n658), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n658), .B1(new_n514), .B2(new_n516), .ZN(new_n931));
  MUX2_X1   g0731(.A(new_n625), .B(new_n621), .S(new_n931), .Z(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT43), .Z(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(KEYINPUT102), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  INV_X1    g0735(.A(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n934), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n663), .ZN(new_n941));
  INV_X1    g0741(.A(new_n923), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n940), .B(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n945));
  XNOR2_X1  g0745(.A(new_n668), .B(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n656), .A2(new_n942), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n655), .A2(new_n649), .A3(new_n923), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT104), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT44), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n656), .A2(new_n952), .A3(new_n953), .A4(new_n942), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n663), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n948), .A2(new_n951), .A3(new_n941), .A4(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT105), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n655), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n653), .A2(new_n654), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n653), .A2(KEYINPUT105), .A3(new_n654), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n662), .A2(KEYINPUT106), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n956), .A2(new_n725), .A3(new_n957), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n946), .B1(new_n969), .B2(new_n725), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n944), .B1(new_n970), .B2(new_n728), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT46), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n765), .B2(new_n442), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n831), .C2(new_n779), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT107), .Z(new_n976));
  OAI21_X1  g0776(.A(new_n372), .B1(new_n486), .B2(new_n752), .ZN(new_n977));
  INV_X1    g0777(.A(new_n774), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G97), .A2(new_n978), .B1(new_n781), .B2(G317), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n833), .B2(new_n827), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n977), .B(new_n980), .C1(G311), .C2(new_n787), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n976), .B(new_n981), .C1(new_n832), .C2(new_n769), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n253), .B1(new_n765), .B2(new_n206), .C1(new_n831), .C2(new_n377), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n774), .A2(new_n213), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n769), .A2(new_n202), .B1(new_n749), .B2(new_n816), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(G150), .C2(new_n771), .ZN(new_n986));
  INV_X1    g0786(.A(G143), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n218), .B2(new_n752), .C1(new_n987), .C2(new_n759), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n982), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n730), .B1(new_n990), .B2(new_n743), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n237), .A2(new_n737), .B1(new_n667), .B2(new_n343), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n744), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(new_n794), .C2(new_n932), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n971), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n725), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n967), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n968), .A2(new_n725), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n668), .B(KEYINPUT113), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n997), .A2(KEYINPUT114), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n653), .A2(new_n794), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n345), .A2(G50), .ZN(new_n1005));
  AOI21_X1  g0805(.A(G45), .B1(new_n1005), .B2(KEYINPUT50), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(KEYINPUT50), .B2(new_n1005), .C1(new_n218), .C2(new_n213), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n241), .A2(G45), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n737), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1010), .B1(new_n227), .B2(new_n253), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(G107), .B2(new_n227), .C1(new_n1012), .C2(new_n666), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT108), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AND3_X1   g0816(.A1(new_n1015), .A2(new_n744), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n761), .A2(G311), .B1(G317), .B2(new_n771), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n787), .A2(G322), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1018), .B(new_n1019), .C1(new_n833), .C2(new_n769), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT110), .Z(new_n1021));
  AOI22_X1  g0821(.A1(new_n1021), .A2(KEYINPUT48), .B1(G294), .B2(new_n766), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n832), .B2(new_n752), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(KEYINPUT48), .B2(new_n1021), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT49), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n781), .A2(G326), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n363), .B1(G116), .B2(new_n978), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT109), .B(G150), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n749), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G77), .A2(new_n766), .B1(new_n771), .B2(G50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n218), .B2(new_n769), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n344), .A2(new_n752), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1036), .A2(new_n372), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G159), .A2(new_n787), .B1(new_n761), .B2(new_n415), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n220), .C2(new_n775), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1031), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT112), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1004), .B(new_n1017), .C1(new_n1042), .C2(new_n743), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1043), .A2(new_n729), .B1(new_n728), .B2(new_n968), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1003), .A2(new_n1044), .ZN(G393));
  INV_X1    g0845(.A(new_n737), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n744), .B1(new_n220), .B2(new_n227), .C1(new_n1046), .C2(new_n248), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n253), .B1(new_n781), .B2(G322), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n442), .B2(new_n752), .C1(new_n779), .C2(new_n769), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n776), .B(new_n1049), .C1(G303), .C2(new_n761), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n787), .A2(G317), .B1(G311), .B2(new_n771), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT52), .Z(new_n1052));
  OAI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(new_n832), .C2(new_n765), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n345), .A2(new_n769), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n787), .A2(G150), .B1(G159), .B2(new_n771), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT51), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n363), .B1(new_n218), .B2(new_n765), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n987), .A2(new_n749), .B1(new_n752), .B2(new_n213), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n824), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n761), .A2(G50), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1053), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n730), .B1(new_n1063), .B2(new_n743), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1047), .B(new_n1064), .C1(new_n923), .C2(new_n794), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n956), .A2(new_n957), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n727), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n969), .A2(new_n1001), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n999), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(G390));
  AND3_X1   g0871(.A1(new_n862), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n886), .A2(new_n860), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n858), .B1(new_n614), .B2(new_n607), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n842), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT39), .B1(new_n1075), .B2(new_n865), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n740), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n253), .B1(new_n752), .B2(new_n377), .ZN(new_n1078));
  INV_X1    g0878(.A(G125), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n827), .A2(new_n822), .B1(new_n749), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n1078), .B(new_n1080), .C1(new_n770), .C2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G128), .A2(new_n787), .B1(new_n761), .B2(G137), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1033), .A2(new_n765), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT53), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G50), .B2(new_n978), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n767), .B1(new_n832), .B2(new_n759), .C1(new_n831), .C2(new_n486), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G97), .A2(new_n770), .B1(new_n781), .B2(G294), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n213), .B2(new_n752), .C1(new_n442), .C2(new_n827), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n1088), .A2(new_n1090), .A3(new_n253), .A4(new_n820), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n743), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n838), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n729), .C1(new_n415), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT116), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1077), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT117), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n875), .B1(new_n806), .B2(new_n894), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n901), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1075), .A2(new_n865), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n802), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n646), .B(new_n1105), .C1(new_n712), .C2(new_n716), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n875), .B1(new_n1106), .B2(new_n894), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1101), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n875), .A2(new_n804), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n706), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n706), .A2(new_n1111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT115), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1103), .A2(new_n1108), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n870), .A2(G330), .A3(new_n804), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n875), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n899), .A2(new_n902), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1104), .A2(new_n1101), .A3(new_n1107), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1099), .B1(new_n728), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n440), .A2(G330), .A3(new_n870), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n906), .A2(new_n616), .A3(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n894), .B(new_n1106), .C1(new_n1117), .C2(new_n1116), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n706), .B2(new_n1111), .ZN(new_n1128));
  AOI211_X1 g0928(.A(KEYINPUT115), .B(new_n1110), .C1(new_n702), .C2(new_n705), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n875), .B1(new_n706), .B2(new_n804), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n896), .B1(new_n1131), .B2(new_n1118), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1126), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1123), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1123), .A2(new_n1133), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1001), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1124), .A2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(new_n1126), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n870), .A2(new_n875), .A3(new_n804), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n862), .B2(new_n865), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n889), .B(G330), .C1(KEYINPUT40), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT118), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n341), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n334), .B2(new_n339), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n320), .A2(new_n857), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1146), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n340), .A2(KEYINPUT118), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n1144), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1148), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1141), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n879), .A2(G330), .A3(new_n889), .A4(new_n1154), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT119), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n905), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n905), .A4(KEYINPUT119), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1138), .A2(new_n1135), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT120), .B1(new_n1162), .B2(KEYINPUT57), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n905), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1159), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1126), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1000), .B1(new_n1169), .B2(KEYINPUT57), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT120), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1172), .C1(new_n1173), .C2(new_n1168), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1163), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1154), .A2(new_n740), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n838), .A2(new_n202), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n372), .B(new_n258), .C1(new_n213), .C2(new_n765), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G58), .A2(new_n978), .B1(new_n781), .B2(G283), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n486), .B2(new_n827), .C1(new_n344), .C2(new_n769), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G68), .C2(new_n753), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n220), .B2(new_n831), .C1(new_n442), .C2(new_n759), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT58), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n759), .A2(new_n1079), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n766), .A2(new_n1081), .B1(new_n770), .B2(G137), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n315), .B2(new_n752), .C1(new_n831), .C2(new_n822), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G128), .C2(new_n771), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT59), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G41), .B1(new_n781), .B2(G124), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G33), .B1(new_n978), .B2(G159), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n370), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G41), .B1(new_n1192), .B2(KEYINPUT3), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1183), .B(new_n1191), .C1(G50), .C2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n730), .B1(new_n1194), .B2(new_n743), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1176), .A2(new_n1177), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1173), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n728), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1175), .A2(new_n1199), .ZN(G375));
  NOR2_X1   g1000(.A1(new_n769), .A2(new_n486), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n827), .A2(new_n832), .B1(new_n749), .B2(new_n833), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G97), .C2(new_n766), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n831), .A2(new_n442), .B1(new_n779), .B2(new_n759), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(new_n1037), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n785), .A2(G77), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n385), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n774), .A2(new_n206), .B1(new_n752), .B2(new_n202), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n372), .B(new_n1208), .C1(G159), .C2(new_n766), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n781), .A2(G128), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G132), .A2(new_n787), .B1(new_n761), .B2(new_n1081), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n770), .A2(G150), .B1(new_n771), .B2(G137), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1214), .A2(new_n746), .B1(G68), .B2(new_n1093), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n730), .B(new_n1215), .C1(new_n1117), .C2(new_n740), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1130), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1132), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1220), .B2(new_n728), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1126), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1133), .A2(new_n946), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G378), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1124), .A2(new_n1136), .A3(KEYINPUT121), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G375), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G384), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1221), .A4(new_n1224), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n971), .A2(new_n1070), .A3(new_n994), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1231), .A2(G396), .A3(G393), .A4(new_n1232), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT122), .Z(G407));
  NAND2_X1  g1034(.A1(new_n1229), .A2(new_n645), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(G409));
  OAI21_X1  g1036(.A(new_n1196), .B1(new_n1167), .B2(new_n727), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1237), .B(new_n1238), .ZN(new_n1239));
  OR3_X1    g1039(.A1(new_n1173), .A2(new_n946), .A3(new_n1168), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1239), .A2(new_n1240), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1175), .A2(G378), .A3(new_n1199), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1175), .A2(new_n1244), .A3(G378), .A4(new_n1199), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1241), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT60), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1133), .B1(new_n1222), .B2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n1001), .C1(new_n1249), .C2(new_n1222), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1221), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1230), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(G384), .A3(new_n1221), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1246), .A2(new_n1248), .A3(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT127), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1241), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1248), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1255), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1257), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1258), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1248), .A2(G2897), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1255), .B(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(new_n1262), .B2(new_n1261), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(KEYINPUT61), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1070), .B1(new_n994), .B2(new_n971), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n798), .B1(new_n1003), .B2(new_n1044), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1275), .A2(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(G390), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(KEYINPUT125), .A4(new_n1232), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1279), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1274), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1264), .B1(new_n1272), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1256), .B2(KEYINPUT63), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1283), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(G405));
  NAND2_X1  g1090(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1243), .A2(new_n1245), .B1(G375), .B2(new_n1291), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1283), .B(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1263), .ZN(G402));
endmodule


