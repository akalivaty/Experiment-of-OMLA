//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n187), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .A4(G128), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT65), .A3(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n192), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT67), .B1(new_n205), .B2(new_n201), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT11), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n208), .B(new_n209), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n203), .B1(KEYINPUT11), .B2(new_n201), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n206), .A2(new_n207), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n216), .A2(KEYINPUT68), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(KEYINPUT68), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n199), .B(new_n204), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n206), .A2(new_n215), .A3(new_n214), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n206), .A2(new_n214), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n207), .A4(new_n215), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(KEYINPUT68), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n195), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n187), .B2(G146), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n189), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n189), .A2(new_n190), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n219), .B(KEYINPUT30), .C1(new_n226), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n226), .B2(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n220), .A2(G131), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n217), .B2(new_n218), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n233), .A2(new_n235), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n219), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n224), .A2(new_n225), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT70), .A3(new_n199), .A4(new_n204), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n239), .A2(new_n244), .A3(new_n246), .A4(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n238), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G116), .B(G119), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n254), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n219), .B(new_n260), .C1(new_n226), .C2(new_n236), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n264), .B(KEYINPUT72), .Z(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n259), .A2(new_n261), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n249), .A2(new_n258), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n241), .A2(new_n243), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n260), .A4(new_n219), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n269), .B1(new_n278), .B2(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT29), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT74), .B(G902), .Z(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n260), .B1(new_n274), .B2(new_n219), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n273), .B2(new_n276), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G472), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n260), .B(new_n238), .C1(new_n250), .C2(new_n249), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n261), .A2(new_n289), .A3(new_n269), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n261), .B2(new_n269), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT31), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n278), .A2(new_n270), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  INV_X1    g110(.A(new_n292), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n259), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n287), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G146), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT16), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT76), .A2(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT76), .A2(G125), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(G140), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G125), .A2(G140), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n307), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n309), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n314), .A2(KEYINPUT16), .A3(G140), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n306), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(KEYINPUT76), .A2(G125), .ZN(new_n317));
  NOR2_X1   g131(.A1(KEYINPUT76), .A2(G125), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n307), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n311), .B1(new_n319), .B2(G140), .ZN(new_n322));
  OAI211_X1 g136(.A(G146), .B(new_n321), .C1(new_n322), .C2(new_n307), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT77), .B(new_n306), .C1(new_n313), .C2(new_n315), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n197), .A3(G119), .ZN(new_n329));
  XNOR2_X1  g143(.A(G119), .B(G128), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n331), .B2(new_n328), .ZN(new_n332));
  INV_X1    g146(.A(G110), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n330), .B(KEYINPUT75), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n338), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n333), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(KEYINPUT78), .ZN(new_n343));
  XOR2_X1   g157(.A(G125), .B(G140), .Z(new_n344));
  OR2_X1    g158(.A1(new_n344), .A2(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(KEYINPUT78), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n343), .A2(new_n323), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT22), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n339), .A2(new_n347), .A3(new_n351), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n282), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT25), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n282), .B2(G234), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n353), .A2(new_n359), .A3(new_n282), .A4(new_n354), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n353), .A2(new_n354), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n358), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT9), .B(G234), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n189), .A2(new_n190), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n192), .B1(new_n370), .B2(new_n198), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G107), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT79), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n372), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n374), .A3(G104), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .A4(new_n373), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n376), .A2(new_n384), .A3(G101), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n371), .A2(new_n378), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n378), .A2(new_n383), .A3(new_n385), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n199), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n241), .A2(new_n389), .A3(KEYINPUT12), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n241), .A2(new_n389), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT12), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n241), .A2(new_n389), .A3(KEYINPUT82), .A4(KEYINPUT12), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n241), .A2(KEYINPUT81), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n247), .A2(new_n399), .A3(new_n240), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT10), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n386), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n388), .A2(KEYINPUT80), .A3(KEYINPUT10), .A4(new_n199), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n379), .A2(new_n381), .A3(new_n373), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n408), .A3(G101), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n407), .A2(new_n235), .A3(new_n233), .A4(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n411));
  INV_X1    g225(.A(new_n199), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n378), .A2(KEYINPUT10), .A3(new_n385), .A4(new_n383), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND4_X1   g228(.A1(new_n403), .A2(new_n404), .A3(new_n410), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n397), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n263), .A2(G227), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n403), .A2(new_n404), .A3(new_n414), .A4(new_n410), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n241), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n401), .B2(new_n415), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n417), .A2(new_n421), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G469), .B1(new_n425), .B2(G902), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n422), .B1(new_n398), .B2(new_n400), .ZN(new_n427));
  INV_X1    g241(.A(new_n423), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n397), .A2(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G469), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n282), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n369), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(G143), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n207), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n187), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  OR3_X1    g254(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n327), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n207), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n437), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n310), .A2(new_n312), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n345), .B1(new_n447), .B2(new_n306), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g263(.A(G113), .B(G122), .Z(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT87), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n372), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n443), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(new_n344), .B2(KEYINPUT19), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n447), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n322), .A2(KEYINPUT86), .A3(KEYINPUT19), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G146), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n323), .B1(new_n438), .B2(new_n440), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n449), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(G475), .A2(G902), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n453), .A2(new_n463), .A3(KEYINPUT88), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n467), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G902), .ZN(new_n473));
  INV_X1    g287(.A(new_n453), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n452), .B1(new_n443), .B2(new_n449), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G122), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G116), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT91), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n481), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(G116), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n481), .A2(new_n480), .B1(new_n484), .B2(KEYINPUT91), .ZN(new_n485));
  OAI21_X1  g299(.A(G107), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G116), .B(G122), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n374), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n197), .A2(G143), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n187), .A2(G128), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n200), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n200), .B1(new_n491), .B2(new_n492), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n486), .B(new_n488), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(KEYINPUT90), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n487), .B(new_n374), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n489), .B(KEYINPUT89), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT13), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n492), .B(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G134), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n491), .A2(new_n503), .A3(new_n200), .A4(new_n492), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(new_n498), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n496), .A2(new_n505), .A3(KEYINPUT92), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n366), .A2(G217), .A3(new_n263), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n510), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n282), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G478), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n511), .A2(new_n282), .A3(new_n513), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n478), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(G234), .A2(G237), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n522), .A2(G952), .A3(new_n263), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n281), .A2(G953), .A3(new_n522), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT21), .B(G898), .Z(new_n527));
  OAI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(G214), .B1(G237), .B2(G902), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT5), .ZN(new_n530));
  INV_X1    g344(.A(G119), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(G116), .ZN(new_n532));
  OAI211_X1 g346(.A(G113), .B(new_n532), .C1(new_n253), .C2(new_n530), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n388), .A2(new_n257), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n407), .A2(new_n258), .A3(new_n409), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT6), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(KEYINPUT83), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n535), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n257), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n387), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT83), .B(new_n539), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(new_n538), .A3(new_n535), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n263), .A2(G224), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT84), .B1(new_n236), .B2(new_n319), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n549));
  AOI211_X1 g363(.A(new_n549), .B(new_n314), .C1(new_n233), .C2(new_n235), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n412), .A2(new_n314), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n549), .B1(new_n243), .B2(new_n314), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n236), .A2(KEYINPUT84), .A3(new_n319), .ZN(new_n555));
  AND4_X1   g369(.A1(new_n552), .A2(new_n554), .A3(new_n555), .A4(new_n547), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n540), .B(new_n546), .C1(new_n553), .C2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n538), .B(KEYINPUT8), .Z(new_n558));
  NAND2_X1  g372(.A1(new_n542), .A2(new_n387), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n534), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n554), .A2(new_n552), .A3(new_n555), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT85), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n562), .A2(KEYINPUT7), .B1(new_n263), .B2(G224), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n562), .B2(KEYINPUT7), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n551), .A2(KEYINPUT7), .A3(new_n552), .A4(new_n547), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n545), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n557), .A2(new_n567), .A3(new_n473), .ZN(new_n568));
  OAI21_X1  g382(.A(G210), .B1(G237), .B2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n557), .A2(new_n567), .A3(new_n473), .A4(new_n569), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n521), .A2(new_n528), .A3(new_n529), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n435), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n305), .A2(new_n365), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(G3));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n300), .B2(new_n282), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n302), .B2(new_n300), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n365), .A3(new_n434), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT93), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n571), .A2(KEYINPUT94), .A3(new_n572), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n529), .B1(new_n571), .B2(KEYINPUT94), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n512), .A2(KEYINPUT95), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n506), .B(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT33), .B1(new_n511), .B2(new_n513), .ZN(new_n590));
  OAI211_X1 g404(.A(G478), .B(new_n282), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT96), .B1(new_n514), .B2(new_n515), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n514), .A2(KEYINPUT96), .A3(new_n515), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n478), .ZN(new_n595));
  INV_X1    g409(.A(new_n528), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n582), .A2(new_n585), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT34), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(new_n372), .ZN(G6));
  INV_X1    g414(.A(new_n468), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT88), .B1(new_n453), .B2(new_n463), .ZN(new_n602));
  INV_X1    g416(.A(new_n467), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n528), .B1(new_n604), .B2(KEYINPUT20), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n520), .A2(new_n469), .A3(new_n477), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT97), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n469), .A2(new_n477), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n596), .B1(new_n610), .B2(new_n471), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .A4(new_n520), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n582), .A2(new_n585), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT35), .B(G107), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT98), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G9));
  NOR2_X1   g431(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n348), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n363), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n361), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT99), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n580), .A2(new_n575), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT37), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n333), .ZN(G12));
  NOR2_X1   g440(.A1(new_n604), .A2(KEYINPUT20), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n523), .B1(new_n525), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n627), .A2(new_n606), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n585), .A2(new_n630), .A3(new_n434), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n305), .A2(new_n623), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XNOR2_X1  g447(.A(new_n629), .B(KEYINPUT39), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n435), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT40), .ZN(new_n636));
  INV_X1    g450(.A(new_n283), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n269), .B1(new_n637), .B2(new_n261), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n259), .B2(new_n298), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n639), .B2(G902), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n303), .B2(new_n304), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n573), .B(KEYINPUT38), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n636), .A2(new_n529), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n520), .ZN(new_n644));
  INV_X1    g458(.A(new_n478), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .A4(new_n623), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n187), .ZN(G45));
  INV_X1    g461(.A(new_n629), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n594), .A2(new_n478), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n585), .A2(new_n649), .A3(new_n434), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n305), .A2(new_n623), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G146), .ZN(G48));
  NAND2_X1  g466(.A1(new_n416), .A2(new_n423), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n421), .B1(new_n397), .B2(new_n424), .ZN(new_n654));
  OAI21_X1  g468(.A(G469), .B1(new_n654), .B2(new_n281), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n433), .A3(KEYINPUT100), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n657), .B(G469), .C1(new_n654), .C2(new_n281), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n369), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n659), .A2(new_n585), .A3(new_n597), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n305), .A3(new_n365), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT101), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT41), .B(G113), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  AND3_X1   g478(.A1(new_n613), .A2(new_n659), .A3(new_n585), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n305), .A3(new_n365), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G116), .ZN(G18));
  NAND2_X1  g481(.A1(new_n656), .A2(new_n658), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n368), .A2(new_n668), .A3(new_n528), .A4(new_n585), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n305), .A2(new_n669), .A3(new_n521), .A4(new_n623), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G119), .ZN(G21));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n284), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n270), .B1(new_n284), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n296), .B1(new_n259), .B2(new_n298), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n294), .B(KEYINPUT103), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n299), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n302), .ZN(new_n681));
  INV_X1    g495(.A(new_n579), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n365), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n478), .A2(new_n684), .A3(new_n520), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n684), .B1(new_n478), .B2(new_n520), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n659), .A3(new_n528), .A4(new_n585), .ZN(new_n688));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n683), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n688), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n579), .B1(new_n680), .B2(new_n302), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n365), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  AND3_X1   g509(.A1(new_n659), .A2(new_n585), .A3(new_n649), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n692), .A3(new_n623), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  OAI21_X1  g512(.A(KEYINPUT107), .B1(new_n303), .B2(new_n304), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n300), .A2(new_n302), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT32), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n699), .A2(new_n704), .A3(new_n287), .ZN(new_n705));
  INV_X1    g519(.A(new_n529), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n573), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n434), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(new_n649), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n365), .A4(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n305), .A2(new_n365), .A3(new_n649), .A4(new_n708), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(KEYINPUT106), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT106), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G131), .ZN(G33));
  AND2_X1   g530(.A1(new_n305), .A2(new_n365), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n630), .A3(new_n708), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(G134), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G36));
  XOR2_X1   g534(.A(new_n425), .B(KEYINPUT45), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(G469), .A2(G902), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n433), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n368), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n634), .ZN(new_n730));
  NOR2_X1   g544(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n645), .A2(new_n594), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n732), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n731), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n682), .A2(new_n700), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n623), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT44), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n730), .A2(new_n742), .A3(new_n707), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  XNOR2_X1  g558(.A(new_n729), .B(KEYINPUT47), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n305), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n365), .A2(new_n595), .A3(new_n629), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n707), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  AOI21_X1  g564(.A(new_n524), .B1(new_n737), .B2(new_n738), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n751), .A2(new_n365), .A3(new_n692), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n707), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n668), .A2(new_n369), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n746), .B2(KEYINPUT114), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n745), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n659), .A2(new_n707), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT117), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n692), .A2(new_n623), .ZN(new_n763));
  INV_X1    g577(.A(new_n641), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n365), .A2(new_n764), .A3(new_n523), .A4(new_n760), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n594), .A2(new_n478), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n762), .A2(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n642), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n752), .A2(new_n706), .A3(new_n768), .A4(new_n659), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT115), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT50), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT116), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(KEYINPUT116), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n758), .B(new_n767), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n718), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n711), .A2(new_n712), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n711), .A2(KEYINPUT106), .A3(new_n712), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n777), .B1(new_n782), .B2(new_n710), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n644), .A2(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n644), .A2(KEYINPUT110), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n627), .B(new_n629), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n305), .A2(new_n608), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n692), .A2(new_n649), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n623), .A3(new_n708), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n670), .A2(new_n661), .A3(new_n666), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n573), .A2(new_n528), .A3(new_n529), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n784), .A2(new_n645), .A3(new_n785), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n595), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n580), .A2(new_n794), .A3(new_n365), .A4(new_n434), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n795), .A2(new_n576), .A3(new_n624), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n694), .A2(new_n790), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n697), .A2(new_n632), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n585), .A2(new_n434), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n621), .A2(new_n629), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n641), .A2(new_n799), .A3(new_n687), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n798), .A2(KEYINPUT52), .A3(new_n651), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n697), .A3(new_n632), .A4(new_n651), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n783), .A2(new_n797), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n623), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n787), .B2(new_n788), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n811), .B2(new_n708), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n715), .A2(new_n718), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n791), .A2(new_n694), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(new_n796), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n689), .A2(new_n693), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n670), .A2(new_n666), .A3(new_n661), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT112), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n813), .A2(new_n806), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n809), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n803), .B(KEYINPUT52), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n808), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n790), .A2(new_n791), .A3(new_n694), .A4(new_n796), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n783), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n806), .B2(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n807), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n821), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT113), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n807), .A2(new_n829), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n807), .A2(new_n829), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n809), .A2(new_n820), .A3(new_n821), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n745), .A2(new_n754), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n775), .B1(new_n839), .B2(new_n753), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n767), .A3(new_n771), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n776), .A2(new_n832), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n705), .A2(new_n365), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n762), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n752), .A2(new_n585), .A3(new_n659), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n765), .A2(new_n478), .A3(new_n594), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n847), .A2(G952), .A3(new_n263), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT118), .Z(new_n850));
  OAI22_X1  g664(.A1(new_n842), .A2(new_n850), .B1(G952), .B2(G953), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n768), .A2(new_n365), .A3(new_n368), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n656), .A2(KEYINPUT49), .A3(new_n658), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT49), .B1(new_n656), .B2(new_n658), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n853), .A2(new_n854), .A3(new_n706), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n764), .A2(new_n852), .A3(new_n734), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n856), .ZN(G75));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n809), .A2(new_n820), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n281), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n860), .B2(new_n569), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n553), .A2(new_n556), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n546), .A2(new_n540), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n557), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT55), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n867), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n282), .B1(new_n809), .B2(new_n820), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(new_n570), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n871), .B2(KEYINPUT119), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n263), .A2(G952), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n871), .B2(KEYINPUT119), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n868), .A2(new_n872), .A3(new_n874), .A4(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(G51));
  NOR2_X1   g693(.A1(new_n860), .A2(new_n722), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT122), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT53), .B1(new_n827), .B2(new_n783), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n806), .A2(new_n819), .A3(new_n796), .A4(new_n815), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n715), .A2(new_n718), .A3(new_n812), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n837), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n859), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n723), .B(KEYINPUT57), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n431), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n873), .B1(new_n881), .B2(new_n892), .ZN(G54));
  AND3_X1   g707(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n601), .A2(new_n602), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n873), .ZN(G60));
  INV_X1    g712(.A(new_n873), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n832), .B2(new_n838), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n589), .A2(new_n590), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n901), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n887), .A2(new_n903), .A3(new_n889), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT60), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n809), .B2(new_n820), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n899), .B1(new_n913), .B2(new_n362), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n619), .B2(new_n913), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g730(.A(new_n263), .B1(new_n527), .B2(G224), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n791), .A2(new_n694), .A3(new_n796), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(new_n263), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n864), .B1(G898), .B2(new_n263), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n920), .B(new_n921), .Z(G69));
  XNOR2_X1  g736(.A(new_n251), .B(new_n458), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n798), .A2(new_n651), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n742), .A2(new_n707), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n843), .A2(new_n585), .A3(new_n687), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(new_n730), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n749), .A2(new_n783), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n263), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n931));
  OR2_X1    g745(.A1(KEYINPUT124), .A2(G900), .ZN(new_n932));
  NAND2_X1  g746(.A1(KEYINPUT124), .A2(G900), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n923), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n646), .A2(new_n924), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n793), .A2(new_n595), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n717), .A2(new_n635), .A3(new_n707), .A4(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n743), .A3(new_n749), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n931), .B1(new_n940), .B2(new_n263), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(new_n923), .ZN(G72));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n940), .B2(new_n919), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n259), .A2(new_n261), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n269), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n270), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT127), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n288), .B2(new_n293), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n944), .B(new_n951), .C1(new_n833), .C2(new_n834), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n944), .B1(new_n929), .B2(new_n919), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n271), .B(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n956), .B2(new_n899), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT126), .B(new_n873), .C1(new_n954), .C2(new_n955), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n948), .B(new_n952), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(G57));
endmodule


