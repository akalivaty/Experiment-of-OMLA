//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n881, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  NAND3_X1  g003(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n212));
  AND4_X1   g011(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n206), .B1(new_n213), .B2(KEYINPUT68), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n209), .A2(new_n211), .A3(new_n207), .A4(new_n212), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n214), .A2(new_n219), .B1(KEYINPUT23), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n220), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n204), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n218), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT70), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n236), .A3(new_n233), .ZN(new_n237));
  INV_X1    g036(.A(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n239));
  AOI21_X1  g038(.A(G190gat), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n235), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n223), .A2(KEYINPUT26), .ZN(new_n245));
  INV_X1    g044(.A(new_n226), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n247), .A3(new_n208), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n217), .A2(new_n218), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n208), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n205), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n249), .A2(new_n250), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n220), .A2(KEYINPUT23), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n255), .A2(new_n204), .A3(new_n228), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G120gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT71), .B(G120gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT72), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n259), .A2(G120gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT1), .B1(new_n267), .B2(new_n260), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(new_n264), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n262), .A2(new_n270), .A3(new_n263), .A4(new_n264), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n229), .A2(new_n258), .A3(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n266), .A2(new_n269), .A3(new_n271), .ZN(new_n274));
  INV_X1    g073(.A(new_n257), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n234), .A2(KEYINPUT70), .B1(new_n240), .B2(KEYINPUT28), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n226), .B1(new_n221), .B2(new_n243), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n276), .A2(new_n237), .B1(new_n277), .B2(new_n245), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(new_n208), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n207), .A2(new_n212), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n209), .A4(new_n211), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n219), .A2(new_n205), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n228), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT25), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n274), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n203), .B1(new_n273), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n272), .B1(new_n229), .B2(new_n258), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n279), .A2(new_n285), .A3(new_n274), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n202), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(new_n293), .B2(KEYINPUT33), .ZN(new_n294));
  XNOR2_X1  g093(.A(G15gat), .B(G43gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G71gat), .ZN(new_n296));
  INV_X1    g095(.A(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n289), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n287), .A2(new_n300), .A3(KEYINPUT32), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n291), .A2(new_n292), .A3(new_n202), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT34), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n202), .B2(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n308), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n291), .A2(new_n292), .A3(new_n202), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n298), .A2(KEYINPUT33), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n305), .A2(new_n314), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n289), .A2(new_n294), .A3(new_n298), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n303), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n315), .B(new_n317), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n313), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G211gat), .B(G218gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  INV_X1    g126(.A(G211gat), .ZN(new_n328));
  INV_X1    g127(.A(G218gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(KEYINPUT22), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n326), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G141gat), .B(G148gat), .Z(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(KEYINPUT2), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n338), .B(new_n337), .C1(new_n342), .C2(KEYINPUT2), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT29), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n333), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT85), .B1(new_n333), .B2(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(G228gat), .ZN(new_n351));
  INV_X1    g150(.A(G233gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n332), .B2(KEYINPUT29), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n341), .A2(new_n343), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n349), .A2(new_n350), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n331), .A2(new_n324), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n331), .A2(new_n324), .ZN(new_n360));
  OR3_X1    g159(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT29), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n361), .B2(new_n344), .ZN(new_n362));
  OAI22_X1  g161(.A1(new_n362), .A2(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n365));
  OAI21_X1  g164(.A(G22gat), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G50gat), .B(G78gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(G106gat), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n369));
  XOR2_X1   g168(.A(new_n368), .B(new_n369), .Z(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n358), .A2(KEYINPUT86), .A3(new_n373), .A4(new_n363), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n366), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n366), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n323), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n229), .B2(new_n258), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n279), .B2(new_n285), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(new_n379), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n332), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(G8gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G36gat), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n333), .B(new_n380), .C1(new_n381), .C2(new_n379), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n387), .B(KEYINPUT79), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n383), .B2(new_n388), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT30), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n272), .A2(new_n356), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n266), .A2(new_n355), .A3(new_n269), .A4(new_n271), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n272), .A2(new_n403), .A3(new_n356), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n344), .B1(new_n341), .B2(new_n343), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n345), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n272), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n272), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n401), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n400), .A2(KEYINPUT82), .A3(new_n402), .A4(new_n404), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n407), .A2(new_n416), .A3(KEYINPUT5), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n399), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n399), .A2(new_n420), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n274), .A2(KEYINPUT4), .A3(new_n355), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n399), .A2(new_n420), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT83), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n401), .A4(new_n414), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT0), .B(G57gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G85gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n429), .A3(new_n434), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n397), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n378), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT35), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n383), .A2(KEYINPUT37), .A3(new_n388), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT37), .B1(new_n383), .B2(new_n388), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT38), .B1(new_n449), .B2(new_n387), .ZN(new_n450));
  INV_X1    g249(.A(new_n448), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n446), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n390), .A2(KEYINPUT38), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n394), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n450), .A2(new_n454), .A3(new_n440), .A4(new_n439), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n427), .A2(new_n414), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n402), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n423), .A2(new_n426), .B1(new_n411), .B2(new_n413), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT87), .B1(new_n459), .B2(new_n401), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT39), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n400), .A2(new_n404), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n401), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n458), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n434), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n396), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(KEYINPUT40), .A3(new_n434), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n436), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n377), .B(new_n455), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n318), .A2(KEYINPUT36), .A3(new_n322), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT36), .B1(new_n318), .B2(new_n322), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n377), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n445), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G113gat), .B(G141gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G169gat), .B(G197gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n485), .B(KEYINPUT12), .Z(new_n486));
  XOR2_X1   g285(.A(G43gat), .B(G50gat), .Z(new_n487));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G29gat), .ZN(new_n490));
  INV_X1    g289(.A(G36gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT14), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n489), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n487), .B2(new_n488), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n488), .B2(new_n487), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n496), .B(KEYINPUT89), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n504), .A2(G1gat), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT16), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n507), .B2(G1gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n506), .B1(new_n505), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(KEYINPUT17), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n503), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n501), .ZN(new_n515));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n516), .B(KEYINPUT90), .Z(new_n517));
  NAND3_X1  g316(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT18), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n518), .A2(KEYINPUT91), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n518), .B2(KEYINPUT91), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n501), .B(new_n511), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n517), .B(KEYINPUT13), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n486), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT18), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n518), .A2(KEYINPUT91), .A3(new_n519), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n525), .A3(new_n529), .A4(new_n486), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G64gat), .ZN(new_n540));
  INV_X1    g339(.A(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G57gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n537), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT97), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  INV_X1    g349(.A(G92gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n552), .A2(new_n553), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n549), .A2(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n550), .A2(new_n551), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n559), .A2(new_n556), .A3(new_n560), .A4(new_n557), .ZN(new_n561));
  INV_X1    g360(.A(new_n553), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n558), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n558), .ZN(new_n565));
  AND4_X1   g364(.A1(new_n559), .A2(new_n556), .A3(new_n560), .A4(new_n557), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n548), .B1(new_n566), .B2(new_n553), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n538), .A2(new_n546), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT10), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n547), .A2(KEYINPUT10), .A3(new_n558), .A4(new_n563), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n571), .A2(new_n572), .B1(G230gat), .B2(G233gat), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n564), .A2(new_n569), .ZN(new_n574));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G120gat), .B(G148gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n225), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G204gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n573), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n575), .B(KEYINPUT98), .Z(new_n583));
  AOI21_X1  g382(.A(new_n583), .B1(new_n571), .B2(new_n572), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n584), .B2(new_n576), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n532), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT96), .ZN(new_n589));
  INV_X1    g388(.A(new_n501), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT93), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n590), .A2(new_n565), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT95), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n503), .A2(new_n565), .A3(new_n512), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n589), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n591), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n588), .A2(KEYINPUT96), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n599), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n514), .B1(KEYINPUT21), .B2(new_n547), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT92), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n611));
  XOR2_X1   g410(.A(G127gat), .B(G155gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G183gat), .B(G211gat), .Z(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n610), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n480), .A2(new_n587), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n441), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G1gat), .ZN(G1324gat));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n621), .A2(new_n396), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(KEYINPUT100), .A3(new_n396), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n627), .A2(new_n626), .A3(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n629), .A2(G8gat), .A3(new_n630), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n635), .A2(KEYINPUT101), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(KEYINPUT101), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n633), .B(new_n634), .C1(new_n636), .C2(new_n637), .ZN(G1325gat));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n474), .B2(new_n475), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n323), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n318), .A2(KEYINPUT36), .A3(new_n322), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(KEYINPUT102), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n621), .A2(G15gat), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(G15gat), .B1(new_n621), .B2(new_n323), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(G1326gat));
  NAND2_X1  g448(.A1(new_n621), .A2(new_n477), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT43), .B(G22gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NAND2_X1  g451(.A1(new_n480), .A2(new_n605), .ZN(new_n653));
  INV_X1    g452(.A(new_n618), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n587), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n490), .A3(new_n623), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659));
  AOI211_X1 g458(.A(KEYINPUT103), .B(new_n377), .C1(new_n397), .C2(new_n441), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n471), .A2(new_n436), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n467), .A2(new_n468), .B1(new_n393), .B2(new_n395), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n477), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n663), .B2(new_n455), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n478), .A2(KEYINPUT103), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n645), .A2(new_n659), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n640), .A3(new_n644), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n442), .A2(new_n668), .A3(new_n477), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n473), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n445), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n605), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n653), .A2(KEYINPUT44), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n655), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(new_n623), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n658), .B1(new_n490), .B2(new_n678), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n656), .A2(new_n491), .A3(new_n396), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT46), .Z(new_n681));
  AND2_X1   g480(.A1(new_n677), .A2(new_n396), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n491), .B2(new_n682), .ZN(G1329gat));
  INV_X1    g482(.A(G43gat), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n656), .A2(new_n684), .A3(new_n323), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n677), .A2(new_n646), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(G43gat), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT47), .B(new_n685), .C1(new_n686), .C2(G43gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n656), .A2(new_n692), .A3(new_n477), .ZN(new_n693));
  INV_X1    g492(.A(new_n655), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n444), .B1(new_n666), .B2(new_n671), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n695), .A2(KEYINPUT44), .A3(new_n606), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n674), .B1(new_n480), .B2(new_n605), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n477), .B(new_n694), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  OAI21_X1  g498(.A(G50gat), .B1(new_n698), .B2(KEYINPUT105), .ZN(new_n700));
  OAI211_X1 g499(.A(KEYINPUT48), .B(new_n693), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n693), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n698), .B2(G50gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(KEYINPUT48), .B2(new_n703), .ZN(G1331gat));
  INV_X1    g503(.A(new_n586), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n526), .A2(new_n531), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n619), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n695), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n623), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n396), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT106), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1333gat));
  INV_X1    g515(.A(new_n709), .ZN(new_n717));
  OAI21_X1  g516(.A(G71gat), .B1(new_n717), .B2(new_n645), .ZN(new_n718));
  INV_X1    g517(.A(G71gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n719), .A3(new_n323), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g521(.A1(new_n709), .A2(new_n477), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n618), .A2(new_n706), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n586), .B(new_n725), .C1(new_n696), .C2(new_n697), .ZN(new_n726));
  INV_X1    g525(.A(new_n623), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n726), .A2(new_n550), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n695), .A2(new_n606), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT51), .Z(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(KEYINPUT107), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n623), .A3(new_n586), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n728), .B1(new_n736), .B2(new_n550), .ZN(G1336gat));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n726), .B2(new_n397), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n729), .B1(new_n675), .B2(new_n676), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT109), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n586), .A4(new_n396), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n741), .A3(G92gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n396), .A2(new_n551), .A3(new_n586), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT108), .Z(new_n744));
  AOI21_X1  g543(.A(KEYINPUT52), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n735), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(G92gat), .B1(new_n726), .B2(new_n397), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(G1337gat));
  NOR3_X1   g550(.A1(new_n726), .A2(new_n297), .A3(new_n645), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n586), .A3(new_n323), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n297), .ZN(G1338gat));
  NOR2_X1   g553(.A1(new_n377), .A2(G106gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n586), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(G106gat), .B1(new_n726), .B2(new_n377), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT53), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n707), .A2(new_n705), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n571), .A2(new_n583), .A3(new_n572), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT54), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n573), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n579), .B1(new_n584), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n571), .A2(new_n572), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n575), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(KEYINPUT110), .A3(KEYINPUT54), .A4(new_n766), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT55), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n768), .A2(new_n773), .A3(new_n776), .A4(new_n770), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT111), .B1(new_n778), .B2(new_n582), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n780), .B(new_n581), .C1(new_n775), .C2(new_n777), .ZN(new_n781));
  INV_X1    g580(.A(new_n485), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n523), .A2(new_n524), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n517), .B1(new_n513), .B2(new_n515), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n530), .A2(new_n785), .ZN(new_n786));
  OR4_X1    g585(.A1(new_n606), .A2(new_n779), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n778), .A2(new_n582), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n780), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n581), .B1(new_n775), .B2(new_n777), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT111), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n706), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n530), .A2(new_n586), .A3(new_n785), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT112), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(KEYINPUT113), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n606), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT113), .B1(new_n792), .B2(new_n794), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n787), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n764), .B1(new_n798), .B2(new_n654), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n378), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n623), .A3(new_n397), .ZN(new_n801));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n532), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n532), .A2(G113gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT114), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n801), .B2(new_n804), .ZN(G1340gat));
  INV_X1    g604(.A(new_n801), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n586), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G120gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n261), .B2(new_n807), .ZN(G1341gat));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n618), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n605), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(G134gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(KEYINPUT116), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n812), .B2(G134gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n812), .A2(new_n817), .A3(G134gat), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI221_X1 g619(.A(new_n815), .B1(new_n813), .B2(new_n816), .C1(new_n818), .C2(new_n820), .ZN(G1343gat));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n654), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n377), .B1(new_n822), .B2(new_n763), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n646), .A2(new_n727), .A3(new_n396), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n706), .A2(new_n790), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n605), .B1(new_n827), .B2(new_n793), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n618), .B1(new_n829), .B2(new_n787), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n477), .B1(new_n830), .B2(new_n764), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT57), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n825), .A2(new_n826), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G141gat), .B1(new_n834), .B2(new_n532), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n823), .A2(new_n623), .A3(new_n645), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n396), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n532), .A2(G141gat), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT117), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g641(.A(G148gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n843), .A3(new_n586), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT59), .B(new_n843), .C1(new_n833), .C2(new_n586), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n477), .A2(new_n824), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n606), .A2(KEYINPUT118), .A3(new_n788), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n605), .B2(new_n790), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n848), .A2(new_n786), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n654), .B1(new_n851), .B2(new_n828), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n852), .B2(new_n763), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n779), .A2(new_n781), .A3(new_n532), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n793), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n606), .A3(new_n795), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n618), .B1(new_n859), .B2(new_n787), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n477), .B1(new_n860), .B2(new_n764), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n853), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n586), .A3(new_n826), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n846), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n844), .B1(new_n845), .B2(new_n864), .ZN(G1345gat));
  INV_X1    g664(.A(new_n837), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n866), .A2(KEYINPUT119), .A3(new_n654), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT119), .B1(new_n866), .B2(new_n654), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n335), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n833), .A2(G155gat), .A3(new_n618), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(G1346gat));
  NOR3_X1   g670(.A1(new_n866), .A2(G162gat), .A3(new_n606), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n873));
  OAI21_X1  g672(.A(G162gat), .B1(new_n834), .B2(new_n606), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT120), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n623), .A2(new_n397), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n800), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n532), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(new_n224), .ZN(G1348gat));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n705), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n225), .ZN(G1349gat));
  NAND2_X1  g681(.A1(new_n238), .A2(new_n239), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n878), .A2(new_n654), .ZN(new_n884));
  MUX2_X1   g683(.A(G183gat), .B(new_n883), .S(new_n884), .Z(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G190gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n878), .A2(new_n606), .ZN(new_n889));
  MUX2_X1   g688(.A(new_n887), .B(new_n888), .S(new_n889), .Z(G1351gat));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n862), .B(KEYINPUT121), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n645), .A2(new_n877), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(new_n532), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n706), .A4(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(G197gat), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n823), .A2(new_n894), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n899), .A2(G197gat), .A3(new_n532), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1352gat));
  NOR3_X1   g700(.A1(new_n899), .A2(G204gat), .A3(new_n705), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906));
  OR3_X1    g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G204gat), .B1(new_n895), .B2(new_n705), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(G1353gat));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT57), .B1(new_n799), .B2(new_n377), .ZN(new_n912));
  INV_X1    g711(.A(new_n853), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n893), .A2(new_n654), .ZN(new_n914));
  AND4_X1   g713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n911), .B1(new_n862), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n919), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n917), .A2(G211gat), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n823), .A2(new_n328), .A3(new_n914), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n862), .A2(new_n911), .A3(new_n914), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n926), .A2(G211gat), .A3(new_n922), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n920), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n923), .A2(new_n929), .A3(KEYINPUT126), .A4(new_n924), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1354gat));
  OAI21_X1  g733(.A(G218gat), .B1(new_n895), .B2(new_n606), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n605), .A2(new_n329), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n899), .B2(new_n936), .ZN(G1355gat));
endmodule


