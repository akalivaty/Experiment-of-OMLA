//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT68), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G137), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n470), .A2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n484), .B1(new_n485), .B2(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT70), .B(G114), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G2105), .ZN(new_n494));
  AND4_X1   g069(.A1(G126), .A2(new_n463), .A3(new_n465), .A4(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G138), .B1(new_n497), .B2(KEYINPUT72), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n482), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n470), .A2(new_n504), .A3(new_n466), .A4(new_n498), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G114), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n492), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(KEYINPUT71), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n496), .A2(new_n501), .A3(new_n505), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n524), .A2(new_n531), .ZN(G166));
  AND2_X1   g107(.A1(new_n529), .A2(G89), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n527), .A2(KEYINPUT73), .A3(new_n528), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  INV_X1    g112(.A(new_n528), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n526), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n539), .A3(G543), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G51), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G168));
  AOI22_X1  g122(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n523), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(KEYINPUT76), .ZN(new_n550));
  INV_X1    g125(.A(new_n540), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(new_n529), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n551), .A2(G52), .B1(new_n553), .B2(G90), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(KEYINPUT76), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  AOI22_X1  g132(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n523), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(G43), .B2(new_n551), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  AND3_X1   g138(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G36), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g144(.A1(new_n518), .A2(new_n520), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  INV_X1    g146(.A(G78), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n570), .A2(new_n571), .B1(new_n572), .B2(new_n517), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI221_X1 g150(.A(KEYINPUT78), .B1(new_n572), .B2(new_n517), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(G651), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n536), .A2(new_n539), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n553), .A2(G91), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  INV_X1    g156(.A(G53), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n540), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  INV_X1    g160(.A(G166), .ZN(G303));
  NAND4_X1  g161(.A1(new_n536), .A2(new_n539), .A3(G49), .A4(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n521), .A2(new_n529), .A3(G87), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  INV_X1    g166(.A(G73), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n570), .A2(new_n591), .B1(new_n592), .B2(new_n517), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n521), .A2(new_n529), .A3(G86), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n529), .A2(G48), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n551), .A2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n553), .A2(G85), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n598), .B(new_n599), .C1(new_n523), .C2(new_n600), .ZN(G290));
  AND3_X1   g176(.A1(new_n521), .A2(G92), .A3(new_n529), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n551), .A2(G54), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n523), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(KEYINPUT79), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(KEYINPUT79), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(G171), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT80), .Z(G284));
  INV_X1    g190(.A(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G299), .A2(new_n611), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n611), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G168), .B2(new_n611), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n610), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g200(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n464), .A2(new_n462), .A3(G2105), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n483), .A2(G135), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n631), .B1(new_n632), .B2(new_n486), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT82), .B(G2096), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2435), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(G14), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT83), .Z(new_n653));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  XOR2_X1   g233(.A(new_n653), .B(KEYINPUT17), .Z(new_n659));
  INV_X1    g234(.A(new_n654), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n659), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  INV_X1    g236(.A(new_n653), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n655), .B1(new_n662), .B2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT85), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2096), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(G227));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT86), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n670), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n676), .B2(new_n672), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n683), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT88), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  XNOR2_X1  g265(.A(KEYINPUT31), .B(G11), .ZN(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G26), .ZN(new_n693));
  INV_X1    g268(.A(new_n486), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G128), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G140), .ZN(new_n696));
  OR2_X1    g271(.A1(G104), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n693), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n693), .B(new_n701), .S(KEYINPUT28), .Z(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G2067), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G19), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n562), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G1341), .Z(new_n707));
  INV_X1    g282(.A(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n692), .B1(new_n708), .B2(G34), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(G34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n480), .B2(new_n692), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2084), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n635), .A2(new_n692), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT97), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(KEYINPUT26), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(KEYINPUT26), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n478), .A2(G105), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n694), .A2(G129), .B1(G141), .B2(new_n483), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n723), .B1(new_n721), .B2(new_n722), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G32), .B(new_n728), .S(G29), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT30), .B(G28), .Z(new_n731));
  OAI22_X1  g306(.A1(new_n729), .A2(new_n730), .B1(G29), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G1961), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n732), .B(new_n735), .C1(G2067), .C2(new_n702), .ZN(new_n736));
  AND4_X1   g311(.A1(new_n703), .A2(new_n717), .A3(new_n719), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G33), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G2105), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G139), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n478), .A2(G103), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT25), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n738), .B1(new_n746), .B2(G29), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G21), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G168), .B2(G16), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n747), .A2(G2072), .B1(G1966), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n692), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n692), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT98), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n750), .B1(G2072), .B2(new_n747), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n692), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n692), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2078), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n749), .A2(G1966), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n704), .A2(KEYINPUT23), .A3(G20), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT23), .ZN(new_n763));
  INV_X1    g338(.A(G20), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G16), .ZN(new_n765));
  INV_X1    g340(.A(G299), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n762), .B(new_n765), .C1(new_n766), .C2(new_n704), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n729), .B2(new_n730), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n754), .A2(new_n755), .B1(G1961), .B2(new_n734), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n737), .A2(new_n761), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G6), .B(G305), .S(G16), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT90), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n773), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n704), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n704), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n783));
  NAND2_X1  g358(.A1(G288), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT91), .A4(new_n589), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n782), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n776), .A2(new_n777), .A3(new_n781), .A4(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G24), .B(G290), .S(G16), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1986), .Z(new_n792));
  OR2_X1    g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n793), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n794));
  INV_X1    g369(.A(G131), .ZN(new_n795));
  INV_X1    g370(.A(G119), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n794), .B1(new_n482), .B2(new_n795), .C1(new_n486), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  INV_X1    g373(.A(G25), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT89), .B1(new_n799), .B2(G29), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n799), .A2(KEYINPUT89), .A3(G29), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT35), .B(G1991), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n802), .B(new_n803), .Z(new_n804));
  NAND3_X1  g379(.A1(new_n790), .A2(new_n792), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT92), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT36), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n776), .A2(new_n781), .A3(new_n789), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n807), .B1(new_n806), .B2(new_n809), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n691), .B(new_n771), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n704), .A2(G4), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n610), .B2(new_n704), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1348), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(G311));
  OR2_X1    g391(.A1(new_n812), .A2(new_n815), .ZN(G150));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n570), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G651), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n553), .A2(G93), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT100), .B(G55), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n822), .B(new_n823), .C1(new_n540), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n562), .A2(new_n825), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n562), .A2(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n610), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n620), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n828), .B1(new_n836), .B2(G860), .ZN(G145));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n838));
  XNOR2_X1  g413(.A(G160), .B(new_n489), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n635), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n728), .B(new_n700), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n501), .A2(new_n505), .A3(new_n513), .A4(new_n512), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n843), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n746), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n844), .A2(new_n746), .A3(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n797), .B(new_n628), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n483), .A2(G142), .ZN(new_n850));
  INV_X1    g425(.A(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n850), .B1(new_n851), .B2(new_n486), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n847), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n847), .B2(new_n848), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n840), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT103), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(new_n840), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n847), .A2(new_n848), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n855), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n847), .A2(new_n848), .A3(new_n856), .ZN(new_n867));
  INV_X1    g442(.A(new_n840), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n864), .B1(new_n863), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n838), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G395));
  NOR2_X1   g451(.A1(new_n825), .A2(G868), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n622), .B(new_n831), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n607), .B(G299), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(KEYINPUT41), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n786), .B(G290), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(KEYINPUT106), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(KEYINPUT106), .ZN(new_n885));
  XOR2_X1   g460(.A(G166), .B(G305), .Z(new_n886));
  OR3_X1    g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n886), .A3(KEYINPUT106), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n881), .B1(new_n878), .B2(new_n882), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n877), .B1(new_n895), .B2(G868), .ZN(G295));
  AOI21_X1  g471(.A(new_n877), .B1(new_n895), .B2(G868), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n898));
  INV_X1    g473(.A(new_n889), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n829), .A2(G286), .A3(new_n830), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G286), .B1(new_n829), .B2(new_n830), .ZN(new_n902));
  OAI21_X1  g477(.A(G301), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n831), .A2(G168), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G171), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n879), .A3(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n903), .A2(new_n905), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n899), .B(new_n906), .C1(new_n907), .C2(new_n882), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n903), .A2(new_n880), .A3(new_n905), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n882), .B1(new_n903), .B2(new_n905), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n889), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n898), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(new_n906), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n889), .B1(new_n915), .B2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n908), .A3(new_n912), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(new_n918), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n908), .A2(new_n911), .A3(new_n912), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n920), .B1(new_n924), .B2(new_n898), .ZN(new_n925));
  AOI211_X1 g500(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n921), .C2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n842), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT110), .B(G40), .Z(new_n932));
  NAND4_X1  g507(.A1(new_n472), .A2(new_n477), .A3(new_n479), .A4(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT111), .Z(new_n937));
  INV_X1    g512(.A(new_n934), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n699), .B(G2067), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(G1996), .B2(new_n728), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n937), .A2(new_n728), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n797), .A2(new_n803), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(G2067), .B2(new_n699), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n934), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n934), .B1(new_n939), .B2(new_n728), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n937), .A2(KEYINPUT46), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n937), .A2(KEYINPUT46), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n941), .B(KEYINPUT112), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n797), .A2(new_n803), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n934), .B1(new_n955), .B2(new_n945), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT48), .Z(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n948), .A2(new_n953), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT127), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n948), .A2(new_n962), .A3(new_n953), .A4(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n842), .A2(KEYINPUT113), .A3(KEYINPUT45), .A4(new_n928), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n515), .A2(new_n928), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n930), .ZN(new_n971));
  INV_X1    g546(.A(G2078), .ZN(new_n972));
  AND4_X1   g547(.A1(new_n477), .A2(new_n472), .A3(new_n479), .A4(new_n932), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n515), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n973), .A3(new_n931), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(KEYINPUT53), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1961), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n515), .B2(new_n928), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n842), .A2(new_n982), .A3(new_n928), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n976), .A2(new_n980), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G171), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT125), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT125), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n990), .A3(G171), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n993));
  INV_X1    g568(.A(G1966), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n978), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n973), .A2(new_n984), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT118), .B(G2084), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n993), .B1(new_n1000), .B2(G286), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n999), .A3(G168), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n993), .B1(new_n1002), .B2(G8), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT62), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G166), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT55), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n933), .B1(new_n970), .B2(new_n930), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1971), .B1(new_n1010), .B2(new_n969), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n983), .A2(new_n985), .A3(G2090), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1009), .B(G8), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n929), .A2(new_n933), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT114), .B1(new_n1014), .B2(new_n1007), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(G8), .C1(new_n929), .C2(new_n933), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n784), .B2(new_n785), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  INV_X1    g599(.A(new_n596), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(G651), .B2(new_n593), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n595), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT115), .B(G86), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n553), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1024), .B(new_n1028), .C1(new_n1031), .C2(new_n1027), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1027), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT49), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1032), .A2(new_n1035), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G288), .A2(new_n1019), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1018), .A2(new_n1038), .A3(new_n1021), .A4(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1013), .A2(new_n1023), .A3(new_n1037), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n933), .B1(KEYINPUT50), .B2(new_n929), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n515), .A2(new_n982), .A3(new_n928), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(KEYINPUT117), .A3(new_n1043), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n755), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1010), .A2(new_n969), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n780), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1009), .B1(new_n1051), .B2(G8), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1041), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1054), .B(new_n1055), .C1(new_n1003), .C2(new_n1001), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n992), .A2(new_n1006), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1038), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1039), .A2(new_n1038), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n1020), .B(new_n1059), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1058), .A2(new_n1060), .A3(new_n1036), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1012), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1007), .B1(new_n1050), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1009), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(G1976), .ZN(new_n1066));
  XOR2_X1   g641(.A(new_n1066), .B(KEYINPUT116), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1028), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1018), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1057), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1009), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1047), .A2(new_n755), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1011), .B1(new_n1072), .B2(new_n1046), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1073), .B2(new_n1007), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1007), .B(G286), .C1(new_n995), .C2(new_n999), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1061), .A3(new_n1013), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1077), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT63), .B1(new_n1063), .B2(new_n1009), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1041), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1075), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1070), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT56), .B(G2072), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1010), .A2(new_n969), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1044), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2067), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1014), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n983), .A2(new_n985), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1094), .B1(new_n1095), .B2(G1348), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n610), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1089), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1089), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n969), .A2(new_n971), .A3(new_n935), .A4(new_n973), .ZN(new_n1107));
  OR2_X1    g682(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1108));
  NAND2_X1  g683(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1108), .B(new_n1109), .C1(new_n929), .C2(new_n933), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n1110), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n562), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1117), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1113), .A2(new_n562), .A3(new_n1119), .A4(new_n1114), .ZN(new_n1120));
  AOI221_X4 g695(.A(KEYINPUT122), .B1(new_n1103), .B2(new_n1106), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n610), .B(KEYINPUT123), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1096), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n834), .A2(KEYINPUT123), .B1(new_n1128), .B2(new_n1096), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1101), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n480), .B(new_n979), .C1(new_n967), .C2(new_n968), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(G40), .A3(new_n931), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n976), .A3(new_n986), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n989), .A2(new_n1137), .A3(new_n991), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1054), .B1(new_n1003), .B2(new_n1001), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1136), .B2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(G171), .B2(new_n987), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(new_n1141), .A3(new_n1053), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1085), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n954), .A2(new_n956), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G290), .B(G1986), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n934), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT126), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n1110), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1119), .B1(new_n1152), .B2(new_n562), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1120), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1124), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1123), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1132), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1101), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1144), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1057), .A2(new_n1064), .A3(new_n1069), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT119), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1084), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT126), .B(new_n1148), .C1(new_n1160), .C2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n964), .B1(new_n1149), .B2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(G401), .A2(G229), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n860), .A2(new_n862), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n1173), .A2(new_n912), .A3(new_n869), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(G319), .ZN(new_n1175));
  NOR3_X1   g749(.A1(new_n1172), .A2(G227), .A3(new_n1175), .ZN(G308));
  OR3_X1    g750(.A1(new_n1172), .A2(G227), .A3(new_n1175), .ZN(G225));
endmodule


