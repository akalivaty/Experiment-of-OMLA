//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n203), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n209), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR4_X1   g0027(.A1(new_n219), .A2(new_n220), .A3(new_n224), .A4(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n222), .A3(G1), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT71), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n223), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT70), .B1(new_n255), .B2(new_n223), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n223), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n223), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n263), .A3(new_n251), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT72), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n258), .A2(new_n263), .A3(KEYINPUT72), .A4(new_n251), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n253), .B1(new_n269), .B2(new_n252), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G58), .A2(G68), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n203), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(G20), .B1(G159), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n222), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT7), .B1(new_n282), .B2(new_n222), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n279), .A2(new_n283), .A3(KEYINPUT77), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(KEYINPUT77), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G68), .ZN(new_n286));
  OAI211_X1 g0086(.A(KEYINPUT16), .B(new_n274), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n261), .A2(new_n262), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT16), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n277), .A2(new_n278), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n202), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n274), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n287), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n270), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(G1), .A3(G13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G274), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  INV_X1    g0104(.A(new_n223), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n299), .ZN(new_n306));
  INV_X1    g0106(.A(new_n302), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(KEYINPUT67), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(G223), .A2(G1698), .ZN(new_n309));
  INV_X1    g0109(.A(G1698), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(G226), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G87), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n311), .A2(new_n282), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n300), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n303), .A2(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n300), .A2(G232), .A3(new_n302), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT78), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n316), .A2(G179), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n316), .B2(new_n318), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n297), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT18), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n297), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n316), .B2(new_n318), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n316), .A2(new_n318), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(G190), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n270), .A2(new_n331), .A3(new_n296), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n270), .A2(new_n331), .A3(KEYINPUT17), .A4(new_n296), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n325), .A2(new_n327), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT73), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n288), .A2(new_n339), .A3(new_n251), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(G68), .C1(G1), .C2(new_n222), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n258), .A2(new_n263), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n222), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n206), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n273), .A2(G50), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n222), .B2(G68), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n343), .B(KEYINPUT11), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n250), .A2(new_n202), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT75), .A2(KEYINPUT12), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n342), .A2(new_n348), .A3(new_n351), .A4(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n230), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G226), .B2(G1698), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n361), .B2(new_n282), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n315), .A2(new_n307), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(new_n315), .B1(new_n363), .B2(G238), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n303), .A2(new_n308), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n368));
  OAI211_X1 g0168(.A(G169), .B(new_n358), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n364), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G179), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n358), .B1(new_n375), .B2(G169), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n357), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n367), .A2(new_n368), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n328), .B1(new_n371), .B2(new_n372), .ZN(new_n380));
  OR3_X1    g0180(.A1(new_n357), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n282), .A2(new_n310), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G238), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n282), .A2(G1698), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G232), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n282), .A2(G107), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n315), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n303), .A2(new_n308), .B1(new_n363), .B2(G244), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n328), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n388), .A2(new_n389), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(G190), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n341), .B(G77), .C1(G1), .C2(new_n222), .ZN(new_n393));
  INV_X1    g0193(.A(new_n252), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT15), .B(G87), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n344), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n397), .A2(new_n289), .B1(new_n206), .B2(new_n250), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n388), .A2(new_n389), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n320), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n388), .A2(new_n389), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n399), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n377), .A2(new_n381), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n336), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n363), .A2(G226), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n366), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n382), .A2(G223), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n282), .A2(G77), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT69), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n384), .B2(G222), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n384), .A2(new_n417), .A3(G222), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n421), .B2(new_n300), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n411), .A2(new_n412), .ZN(new_n423));
  OAI21_X1  g0223(.A(G200), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n420), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n415), .B(new_n414), .C1(new_n425), .C2(new_n418), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n315), .B1(new_n412), .B2(new_n411), .ZN(new_n427));
  INV_X1    g0227(.A(new_n423), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(G190), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n269), .A2(G50), .ZN(new_n431));
  INV_X1    g0231(.A(new_n344), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n394), .A2(new_n432), .B1(G150), .B2(new_n273), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n205), .B2(new_n222), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n343), .B1(new_n242), .B2(new_n250), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT9), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(KEYINPUT9), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n430), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT74), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT10), .B1(new_n430), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI221_X1 g0243(.A(new_n430), .B1(new_n441), .B2(KEYINPUT10), .C1(new_n438), .C2(new_n439), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n320), .B1(new_n422), .B2(new_n423), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n427), .A2(new_n404), .A3(new_n428), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n436), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n409), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n451));
  OAI211_X1 g0251(.A(G250), .B(new_n310), .C1(new_n280), .C2(new_n281), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G294), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n455), .A2(new_n457), .B1(new_n305), .B2(new_n299), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n454), .A2(new_n315), .B1(new_n458), .B2(G264), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n268), .A2(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n306), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(G179), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n320), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n313), .A2(G20), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n280), .B2(new_n281), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n222), .A2(G87), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n275), .B2(new_n276), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT22), .B1(new_n475), .B2(KEYINPUT84), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n469), .B(KEYINPUT84), .C1(new_n281), .C2(new_n280), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n470), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n477), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n472), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G107), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT23), .A3(G20), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT23), .B1(new_n485), .B2(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n487), .A2(new_n488), .B1(G20), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT24), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n472), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n470), .A2(new_n481), .ZN(new_n493));
  AND4_X1   g0293(.A1(KEYINPUT85), .A2(new_n493), .A3(KEYINPUT22), .A4(new_n477), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT85), .B1(new_n482), .B2(new_n477), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  INV_X1    g0297(.A(new_n490), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n288), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n268), .A2(G33), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n258), .A2(new_n263), .A3(new_n251), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n485), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n250), .A2(new_n485), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT25), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n468), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n484), .A2(KEYINPUT24), .A3(new_n490), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n289), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n466), .A2(new_n328), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G190), .B2(new_n466), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G97), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n502), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  AND2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n485), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n273), .A2(G77), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n485), .B1(new_n291), .B2(new_n292), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n289), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n250), .A2(new_n517), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n518), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n310), .C1(new_n280), .C2(new_n281), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n275), .A2(new_n276), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(KEYINPUT4), .A3(G244), .A4(new_n310), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n534), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n315), .ZN(new_n540));
  INV_X1    g0340(.A(new_n463), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n457), .B1(new_n541), .B2(new_n461), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(G257), .A3(new_n300), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n465), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n320), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n544), .B1(new_n539), .B2(new_n315), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n404), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n531), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(G200), .ZN(new_n551));
  OAI21_X1  g0351(.A(G107), .B1(new_n279), .B2(new_n283), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n524), .A2(G20), .B1(G77), .B2(new_n273), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(new_n289), .B1(new_n517), .B2(new_n250), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(G190), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n551), .A2(new_n518), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n255), .A2(new_n223), .B1(G20), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n537), .B(new_n222), .C1(G33), .C2(new_n517), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT20), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(G116), .B2(new_n251), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n501), .A2(G116), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n341), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n458), .A2(G270), .B1(new_n306), .B2(new_n464), .ZN(new_n569));
  OAI211_X1 g0369(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n570));
  OAI211_X1 g0370(.A(G257), .B(new_n310), .C1(new_n280), .C2(new_n281), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n315), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G169), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n559), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(G200), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n574), .A3(G190), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n568), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n569), .A2(G179), .A3(new_n574), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n566), .B1(new_n338), .B2(new_n340), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n565), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n320), .B1(new_n569), .B2(new_n574), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(KEYINPUT21), .C1(new_n582), .C2(new_n565), .ZN(new_n585));
  AND4_X1   g0385(.A1(new_n577), .A2(new_n580), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n344), .B2(new_n517), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n222), .A2(G68), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n282), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n222), .B1(new_n359), .B2(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n521), .A2(new_n313), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n590), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n396), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n597), .A2(new_n288), .B1(new_n251), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n502), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT83), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(G87), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT83), .B1(new_n502), .B2(new_n313), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g0404(.A1(G238), .A2(G1698), .ZN(new_n605));
  INV_X1    g0405(.A(G244), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G1698), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n280), .C2(new_n281), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n489), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT80), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT80), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n611), .A3(new_n489), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n315), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n300), .A2(G274), .A3(new_n457), .ZN(new_n614));
  AND2_X1   g0414(.A1(G33), .A2(G41), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n460), .B(G250), .C1(new_n615), .C2(new_n223), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT79), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT79), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n614), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n613), .A2(new_n621), .A3(new_n378), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n300), .B1(new_n609), .B2(KEYINPUT80), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(new_n612), .B1(new_n618), .B2(new_n620), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(G200), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n604), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n613), .A2(new_n621), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n404), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n320), .B1(new_n613), .B2(new_n621), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT81), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(G169), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(G179), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT81), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n502), .A2(new_n396), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n599), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n630), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n558), .A2(new_n586), .A3(new_n626), .A4(new_n637), .ZN(new_n638));
  NOR4_X1   g0438(.A1(new_n450), .A2(new_n509), .A3(new_n516), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n447), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n443), .A2(new_n444), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n334), .A2(new_n335), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n357), .A2(new_n379), .A3(new_n380), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n377), .B2(new_n407), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI211_X1 g0445(.A(KEYINPUT18), .B(new_n322), .C1(new_n270), .C2(new_n296), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n326), .B1(new_n297), .B2(new_n323), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n640), .B1(new_n641), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n531), .A2(new_n547), .A3(new_n549), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n637), .A2(new_n651), .A3(new_n626), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n631), .A2(new_n632), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n636), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n604), .A2(new_n625), .B1(new_n654), .B2(new_n636), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n651), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n515), .A2(new_n558), .A3(new_n656), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n577), .A2(new_n583), .A3(new_n585), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n512), .A2(new_n506), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n468), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT87), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n508), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n550), .A2(new_n557), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n491), .A2(new_n499), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n507), .B1(new_n668), .B2(new_n289), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n669), .B2(new_n514), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n666), .A2(new_n670), .A3(new_n671), .A4(new_n656), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n659), .B1(new_n664), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n650), .B1(new_n450), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT88), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n268), .A2(new_n222), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n568), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n661), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n577), .A2(new_n580), .A3(new_n583), .A4(new_n585), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n684), .B(G330), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n687), .A2(new_n686), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(KEYINPUT90), .A3(G330), .A4(new_n684), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n681), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n509), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n515), .B(new_n508), .C1(new_n669), .C2(new_n681), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n509), .A2(new_n681), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n515), .A2(new_n508), .A3(new_n681), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(new_n665), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n592), .A2(G116), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT91), .Z(new_n704));
  INV_X1    g0504(.A(new_n225), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n221), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n652), .A2(KEYINPUT94), .A3(new_n657), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n626), .A4(new_n655), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n656), .A2(KEYINPUT93), .A3(KEYINPUT26), .A4(new_n651), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT94), .B1(new_n652), .B2(new_n657), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n712), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n655), .B1(new_n660), .B2(new_n663), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n681), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n664), .A2(new_n672), .ZN(new_n722));
  INV_X1    g0522(.A(new_n659), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n694), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n721), .B1(KEYINPUT29), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n546), .A2(new_n466), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n608), .A2(new_n611), .A3(new_n489), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n611), .B1(new_n608), .B2(new_n489), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n728), .A2(new_n729), .A3(new_n300), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n614), .A2(new_n619), .A3(new_n616), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n619), .B1(new_n614), .B2(new_n616), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n404), .B(new_n575), .C1(new_n730), .C2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n726), .B1(new_n727), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n581), .A2(new_n624), .A3(new_n548), .A4(new_n459), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n613), .A2(new_n621), .A3(new_n459), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .A3(new_n581), .A4(new_n548), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n540), .A2(new_n545), .B1(new_n459), .B2(new_n465), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n613), .B2(new_n621), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n741), .A2(KEYINPUT92), .A3(new_n575), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n735), .A2(new_n738), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n694), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n738), .A2(new_n740), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n727), .A2(new_n734), .ZN(new_n749));
  OAI211_X1 g0549(.A(KEYINPUT31), .B(new_n694), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n747), .B(new_n750), .C1(new_n700), .C2(new_n638), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n725), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n710), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n249), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n268), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n706), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(G330), .B1(new_n691), .B2(new_n684), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n761), .B1(new_n693), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(G20), .B(new_n765), .C1(new_n691), .C2(new_n684), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n705), .A2(new_n282), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n767), .A2(G355), .B1(new_n560), .B2(new_n705), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n247), .A2(new_n456), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n705), .A2(new_n535), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G45), .B2(new_n221), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n765), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n223), .B1(G20), .B2(new_n320), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n222), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(G303), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n282), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT96), .Z(new_n781));
  NAND2_X1  g0581(.A1(G20), .A2(G179), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n378), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(G190), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G200), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G311), .A2(new_n785), .B1(new_n787), .B2(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n328), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n378), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n222), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n789), .A2(G326), .B1(G294), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n784), .A2(new_n328), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n781), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n777), .A2(new_n378), .A3(new_n328), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT97), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n777), .A2(new_n378), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n802), .A2(G329), .B1(G283), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT98), .ZN(new_n806));
  INV_X1    g0606(.A(new_n798), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G159), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n803), .A2(new_n485), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n791), .A2(new_n517), .B1(new_n778), .B2(new_n313), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n809), .A2(new_n282), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n789), .ZN(new_n813));
  INV_X1    g0613(.A(new_n787), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n242), .A2(new_n813), .B1(new_n814), .B2(new_n201), .ZN(new_n815));
  INV_X1    g0615(.A(new_n795), .ZN(new_n816));
  INV_X1    g0616(.A(new_n785), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n202), .A2(new_n816), .B1(new_n817), .B2(new_n206), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n797), .A2(new_n806), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n774), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n776), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n760), .B1(new_n766), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n763), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT99), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n722), .A2(new_n723), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n406), .A2(new_n681), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n681), .B1(new_n393), .B2(new_n398), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n392), .B2(new_n400), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n829), .B2(new_n406), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(new_n681), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n673), .B2(new_n694), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n753), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT100), .Z(new_n836));
  AOI21_X1  g0636(.A(new_n760), .B1(new_n834), .B2(new_n753), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n774), .A2(new_n764), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n761), .B1(new_n206), .B2(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n560), .A2(new_n817), .B1(new_n813), .B2(new_n779), .ZN(new_n841));
  INV_X1    g0641(.A(G283), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n842), .A2(new_n816), .B1(new_n814), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n803), .A2(new_n313), .ZN(new_n845));
  INV_X1    g0645(.A(new_n778), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G107), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n535), .B1(new_n792), .B2(G97), .ZN(new_n848));
  INV_X1    g0648(.A(G311), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n847), .B(new_n848), .C1(new_n801), .C2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n841), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n787), .B1(new_n785), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(G137), .ZN(new_n853));
  INV_X1    g0653(.A(G150), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n853), .B2(new_n813), .C1(new_n854), .C2(new_n816), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n535), .B1(new_n778), .B2(new_n242), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n791), .A2(new_n201), .B1(new_n803), .B2(new_n202), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n802), .C2(G132), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n851), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n840), .B1(new_n860), .B2(new_n821), .C1(new_n831), .C2(new_n765), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n838), .A2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n757), .A2(new_n268), .ZN(new_n863));
  INV_X1    g0663(.A(G330), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n747), .B(new_n865), .C1(new_n700), .C2(new_n638), .ZN(new_n866));
  OAI21_X1  g0666(.A(G169), .B1(new_n367), .B2(new_n368), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(KEYINPUT76), .A3(KEYINPUT14), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n373), .A3(new_n369), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n357), .B(new_n694), .C1(new_n869), .C2(new_n643), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n357), .A2(new_n694), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n377), .A2(new_n381), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n830), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n274), .B1(new_n284), .B2(new_n286), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n290), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n343), .A3(new_n287), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n679), .B1(new_n270), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n336), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n297), .A2(new_n680), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n324), .A2(new_n880), .A3(new_n881), .A4(new_n332), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n270), .A2(new_n331), .A3(new_n296), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n322), .B1(new_n270), .B2(new_n877), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n883), .A2(new_n884), .A3(new_n878), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n880), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n336), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n324), .A2(new_n880), .A3(new_n332), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n882), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n874), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n866), .A2(new_n873), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT103), .B1(new_n866), .B2(new_n873), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n883), .A2(new_n878), .ZN(new_n901));
  INV_X1    g0701(.A(new_n884), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n881), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n882), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n878), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n648), .B2(new_n642), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n900), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n879), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n894), .A2(KEYINPUT40), .B1(new_n899), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT104), .Z(new_n912));
  INV_X1    g0712(.A(new_n866), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n450), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n864), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n912), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT102), .ZN(new_n917));
  INV_X1    g0717(.A(new_n827), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n724), .B2(new_n831), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n870), .A2(new_n872), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n673), .A2(new_n694), .A3(new_n830), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT102), .B(new_n920), .C1(new_n923), .C2(new_n918), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n924), .A3(new_n910), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n887), .B2(new_n893), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n908), .A2(KEYINPUT39), .A3(new_n909), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n869), .A2(new_n357), .A3(new_n681), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n679), .B1(new_n646), .B2(new_n647), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n721), .B(new_n449), .C1(KEYINPUT29), .C2(new_n724), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n650), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n863), .B1(new_n916), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n916), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n223), .A2(new_n222), .A3(new_n560), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n524), .B(KEYINPUT101), .Z(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT35), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n942), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  NAND2_X1  g0746(.A1(new_n271), .A2(G77), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n243), .B1(new_n221), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(G1), .A3(new_n249), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n939), .A2(new_n946), .A3(new_n949), .ZN(G367));
  NAND2_X1  g0750(.A1(new_n531), .A2(new_n694), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n558), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n651), .A2(new_n694), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n701), .A2(new_n699), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT106), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n955), .A2(new_n957), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n954), .B1(new_n701), .B2(new_n699), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT44), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n962), .B(new_n954), .C1(new_n701), .C2(new_n699), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n958), .A2(new_n959), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(KEYINPUT108), .A3(new_n698), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n960), .B(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n698), .A2(KEYINPUT108), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n955), .B(new_n957), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT108), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n693), .A2(new_n969), .A3(new_n697), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT107), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n665), .A2(new_n694), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n701), .B1(new_n697), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n973), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n754), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n706), .B(KEYINPUT41), .Z(new_n978));
  OAI21_X1  g0778(.A(new_n758), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n954), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n701), .A2(KEYINPUT42), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n550), .B1(new_n952), .B2(new_n508), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n681), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT42), .B1(new_n701), .B2(new_n980), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n604), .A2(new_n681), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n655), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n656), .B2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n989), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n989), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n985), .A2(new_n993), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n698), .A2(new_n980), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n979), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n237), .A2(new_n770), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n775), .B1(new_n225), .B2(new_n396), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n760), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n789), .A2(G143), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n817), .B2(new_n242), .C1(new_n854), .C2(new_n814), .ZN(new_n1003));
  INV_X1    g0803(.A(G159), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n816), .A2(new_n1004), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n535), .B1(new_n798), .B2(new_n853), .C1(new_n206), .C2(new_n803), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n792), .A2(G68), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n201), .B2(new_n778), .ZN(new_n1008));
  NOR4_X1   g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT111), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT46), .B1(new_n846), .B2(G116), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT110), .B(G317), .Z(new_n1012));
  OAI221_X1 g0812(.A(new_n282), .B1(new_n803), .B2(new_n517), .C1(new_n798), .C2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(G107), .C2(new_n792), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G294), .A2(new_n795), .B1(new_n789), .B2(G311), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G283), .A2(new_n785), .B1(new_n787), .B2(G303), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n846), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT109), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1010), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT47), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1001), .B1(new_n1021), .B2(new_n774), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n773), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n998), .A2(new_n1024), .ZN(G387));
  NAND3_X1  g0825(.A1(new_n695), .A2(new_n696), .A3(new_n773), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n770), .B1(new_n233), .B2(new_n456), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n767), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1027), .B1(new_n704), .B2(new_n1028), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n252), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT50), .B1(new_n252), .B2(G50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n704), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1029), .A2(new_n1033), .B1(new_n485), .B2(new_n705), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n775), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n760), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n242), .A2(new_n814), .B1(new_n813), .B2(new_n1004), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n394), .B2(new_n795), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n535), .B1(new_n798), .B2(new_n854), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n846), .A2(G77), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n396), .B2(new_n791), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(G97), .C2(new_n804), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1038), .B(new_n1042), .C1(new_n202), .C2(new_n817), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n535), .B1(new_n807), .B2(G326), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n791), .A2(new_n842), .B1(new_n778), .B2(new_n843), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G303), .A2(new_n785), .B1(new_n795), .B2(G311), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n789), .A2(G322), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n814), .C2(new_n1012), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1044), .B1(new_n560), .B2(new_n803), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1043), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n774), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n976), .A2(new_n759), .B1(new_n1026), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n755), .A2(new_n976), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n706), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n755), .A2(new_n976), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n965), .A3(new_n971), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n972), .A2(new_n755), .A3(new_n976), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n1063), .A3(new_n706), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n980), .A2(new_n773), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n770), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n775), .B1(new_n517), .B2(new_n225), .C1(new_n241), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n760), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G311), .A2(new_n787), .B1(new_n789), .B2(G317), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT52), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n535), .B(new_n810), .C1(G322), .C2(new_n807), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n792), .A2(G116), .B1(new_n846), .B2(G283), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n843), .B2(new_n817), .C1(new_n779), .C2(new_n816), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n282), .B(new_n845), .C1(G143), .C2(new_n807), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n792), .A2(G77), .B1(new_n846), .B2(G68), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n242), .B2(new_n816), .C1(new_n252), .C2(new_n817), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G150), .A2(new_n789), .B1(new_n787), .B2(G159), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT51), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1070), .A2(new_n1074), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1068), .B1(new_n1081), .B2(new_n774), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n972), .A2(new_n759), .B1(new_n1065), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1064), .A2(new_n1083), .ZN(G390));
  NOR2_X1   g0884(.A1(new_n913), .A2(new_n864), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n873), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n920), .B1(new_n923), .B2(new_n918), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1088), .A2(new_n929), .B1(new_n927), .B2(new_n928), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n336), .A2(new_n888), .B1(new_n891), .B2(new_n882), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n909), .B1(new_n1090), .B2(KEYINPUT38), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n929), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n829), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n407), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n681), .B(new_n1094), .C1(new_n719), .C2(new_n720), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n827), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1092), .B1(new_n1096), .B2(new_n920), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n920), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1091), .A2(new_n929), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n751), .A2(G330), .A3(new_n831), .A4(new_n920), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n832), .A2(new_n827), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n930), .B1(new_n1103), .B2(new_n920), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n927), .A2(new_n928), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1101), .B(new_n1102), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n449), .A2(new_n1085), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n935), .A2(new_n650), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT112), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n866), .A2(new_n1111), .A3(G330), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n831), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n866), .B2(G330), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n921), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT113), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1095), .A2(new_n827), .A3(new_n1102), .ZN(new_n1118));
  OAI211_X1 g0918(.A(KEYINPUT113), .B(new_n921), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n920), .B1(new_n752), .B2(new_n831), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1103), .B1(new_n1087), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1110), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1108), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1098), .A2(new_n1123), .A3(new_n1107), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n706), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1098), .A2(new_n759), .A3(new_n1107), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n839), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n760), .B1(new_n394), .B2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT114), .Z(new_n1131));
  NAND2_X1  g0931(.A1(new_n846), .A2(G150), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G125), .B2(new_n802), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n787), .A2(G132), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT115), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n789), .B1(new_n785), .B2(new_n1137), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n535), .B1(new_n803), .B2(new_n242), .C1(new_n791), .C2(new_n1004), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G137), .B2(new_n795), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n282), .B1(new_n803), .B2(new_n202), .C1(new_n313), .C2(new_n778), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n802), .B2(G294), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G107), .A2(new_n795), .B1(new_n789), .B2(G283), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n517), .C2(new_n817), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n787), .A2(G116), .B1(G77), .B2(new_n792), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT116), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1141), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n821), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT118), .Z(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1106), .B2(new_n765), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1128), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1127), .A2(new_n1155), .ZN(G378));
  XNOR2_X1  g0956(.A(new_n1110), .B(KEYINPUT121), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1126), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n448), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n443), .A2(new_n444), .A3(new_n447), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n679), .B1(new_n431), .B2(new_n435), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT119), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1160), .A2(new_n1165), .A3(new_n1162), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n911), .B2(new_n864), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n899), .A2(new_n910), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT40), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1091), .B2(new_n874), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1171), .B(G330), .C1(new_n1172), .C2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n934), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1170), .A2(new_n925), .A3(new_n1175), .A4(new_n933), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(KEYINPUT57), .A3(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n706), .B1(new_n1158), .B2(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1126), .A2(new_n1157), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n759), .A3(new_n1178), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n760), .B1(G50), .B2(new_n1129), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n535), .A2(G41), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n242), .B1(G33), .B2(G41), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n804), .A2(G58), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1007), .A2(new_n1040), .A3(new_n1186), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G283), .B2(new_n802), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G97), .A2(new_n795), .B1(new_n789), .B2(G116), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G107), .A2(new_n787), .B1(new_n785), .B2(new_n598), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n789), .A2(G125), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G128), .A2(new_n787), .B1(new_n785), .B2(G137), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1137), .A2(new_n846), .B1(G150), .B2(new_n792), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n795), .A2(G132), .ZN(new_n1200));
  AND4_X1   g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n804), .A2(G159), .ZN(new_n1204));
  AOI211_X1 g1004(.A(G33), .B(G41), .C1(new_n807), .C2(G124), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1208), .B2(new_n774), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1169), .B2(new_n765), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT120), .B1(new_n1184), .B2(new_n1210), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1180), .A2(new_n1183), .B1(new_n1211), .B2(new_n1212), .ZN(G375));
  INV_X1    g1013(.A(new_n978), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1120), .A2(new_n1122), .A3(new_n1110), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1124), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n758), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n921), .A2(new_n764), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n760), .B1(G68), .B2(new_n1129), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n485), .A2(new_n817), .B1(new_n816), .B2(new_n560), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n842), .A2(new_n814), .B1(new_n813), .B2(new_n843), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n792), .A2(new_n598), .B1(new_n846), .B2(G97), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n535), .B1(new_n804), .B2(G77), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n801), .C2(new_n779), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  AOI22_X1  g1026(.A1(G132), .A2(new_n789), .B1(new_n795), .B2(new_n1137), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n853), .B2(new_n814), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT123), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n802), .A2(G128), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n785), .A2(G150), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n282), .B1(new_n804), .B2(G58), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n792), .A2(G50), .B1(new_n846), .B2(G159), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1229), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1219), .B1(new_n1235), .B2(new_n774), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1217), .B1(new_n1218), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1216), .A2(new_n1237), .ZN(G381));
  NAND2_X1  g1038(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1179), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n707), .B1(new_n1242), .B2(new_n1182), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1184), .A2(new_n1210), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT120), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1184), .A2(KEYINPUT120), .A3(new_n1210), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1241), .A2(new_n1243), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1127), .A2(new_n1155), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OR2_X1    g1050(.A1(G393), .A2(G396), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n1251), .A2(G384), .A3(G390), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G387), .A2(new_n1250), .A3(G381), .A4(new_n1252), .ZN(G407));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  INV_X1    g1054(.A(new_n1244), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1181), .A2(new_n1214), .A3(new_n1182), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1249), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(G375), .B2(new_n1249), .ZN(new_n1259));
  INV_X1    g1059(.A(G343), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(G213), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1215), .B1(new_n1123), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(KEYINPUT124), .B(new_n1215), .C1(new_n1123), .C2(new_n1262), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1215), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n707), .B1(new_n1267), .B2(KEYINPUT60), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(G384), .A3(new_n1237), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1269), .B2(new_n1237), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1259), .A2(new_n1261), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(KEYINPUT62), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1259), .A2(new_n1272), .A3(new_n1276), .A4(new_n1261), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1261), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(G2897), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1269), .A2(new_n1237), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1269), .A2(G384), .A3(new_n1237), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1279), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(G378), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1248), .B2(G378), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1289), .B2(new_n1278), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G393), .A2(G396), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1251), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT126), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1251), .A2(new_n1295), .A3(new_n1292), .ZN(new_n1296));
  INV_X1    g1096(.A(G390), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(G387), .A2(new_n1297), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n979), .A2(new_n997), .B1(new_n1023), .B2(new_n1022), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1299), .A2(G390), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1294), .B(new_n1296), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G387), .A2(KEYINPUT127), .A3(new_n1297), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1299), .B2(G390), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(G390), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(new_n1304), .A3(new_n1305), .A4(new_n1293), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1301), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1291), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1273), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1287), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1280), .A2(new_n1286), .A3(KEYINPUT125), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1273), .A2(new_n1309), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1307), .A2(KEYINPUT61), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1310), .A2(new_n1315), .A3(new_n1316), .A4(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1318), .ZN(G405));
  NOR2_X1   g1119(.A1(G375), .A2(new_n1249), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1248), .A2(G378), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1307), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1320), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1301), .A2(new_n1306), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1322), .A2(new_n1272), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1272), .B1(new_n1322), .B2(new_n1325), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


