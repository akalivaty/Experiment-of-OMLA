//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(new_n202), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(KEYINPUT65), .A2(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(KEYINPUT65), .A2(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G58), .B2(G232), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G107), .A2(G264), .ZN(new_n227));
  NAND4_X1  g0027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G97), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n253), .B(new_n254), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G238), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n262), .A3(G274), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT74), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  INV_X1    g0074(.A(new_n215), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(new_n261), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT74), .B1(new_n276), .B2(new_n270), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n267), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT13), .B1(new_n260), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT75), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n258), .A2(new_n259), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n273), .A2(new_n277), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n267), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(KEYINPUT75), .B(KEYINPUT13), .C1(new_n260), .C2(new_n278), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G169), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n285), .A2(new_n286), .A3(new_n289), .A4(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n279), .A2(G179), .A3(new_n284), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT67), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n296));
  AND4_X1   g0096(.A1(KEYINPUT68), .A2(new_n294), .A3(new_n215), .A4(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n293), .A2(KEYINPUT67), .B1(G1), .B2(G13), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT68), .B1(new_n298), .B2(new_n296), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n216), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n221), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n302), .B1(new_n303), .B2(new_n304), .C1(new_n305), .C2(new_n216), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g0107(.A(new_n307), .B(KEYINPUT11), .Z(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(new_n216), .A3(G1), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n294), .A2(new_n215), .A3(new_n296), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n298), .A2(KEYINPUT68), .A3(new_n296), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n263), .A2(G20), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(G68), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT77), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT12), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g0122(.A(new_n310), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT12), .B1(new_n305), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n317), .A2(new_n318), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n318), .B1(new_n317), .B2(new_n326), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n308), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n292), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n279), .A2(G190), .A3(new_n284), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n285), .A2(G200), .A3(new_n286), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n335));
  INV_X1    g0135(.A(G107), .ZN(new_n336));
  INV_X1    g0136(.A(G232), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n335), .B1(new_n336), .B2(new_n252), .C1(new_n256), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n259), .ZN(new_n339));
  INV_X1    g0139(.A(G244), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n271), .B1(new_n265), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n338), .B2(new_n259), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G20), .A2(G77), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT8), .B(G58), .ZN(new_n351));
  INV_X1    g0151(.A(new_n301), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n350), .B1(new_n351), .B2(new_n352), .C1(new_n304), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n310), .A2(new_n303), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT70), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n355), .A2(KEYINPUT70), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n300), .A2(new_n354), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n315), .A2(G77), .A3(new_n316), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n349), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n343), .A2(G200), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n346), .A2(G190), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n362), .A2(new_n359), .A3(new_n358), .A4(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n331), .A2(new_n334), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n252), .A2(G222), .A3(new_n255), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n252), .A2(G223), .A3(G1698), .ZN(new_n368));
  AND2_X1   g0168(.A1(KEYINPUT3), .A2(G33), .ZN(new_n369));
  NOR2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G77), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n259), .ZN(new_n374));
  INV_X1    g0174(.A(new_n271), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(G226), .B2(new_n266), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(G179), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n203), .A2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n301), .A2(G150), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT69), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n351), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  OR3_X1    g0183(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT8), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n379), .B(new_n380), .C1(new_n385), .C2(new_n304), .ZN(new_n386));
  INV_X1    g0186(.A(G50), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(new_n300), .B1(new_n387), .B2(new_n310), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n315), .A2(G50), .A3(new_n316), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n378), .B(new_n391), .C1(new_n344), .C2(new_n377), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n374), .A2(G190), .A3(new_n376), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT71), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT71), .A4(G190), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT9), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n388), .A2(new_n399), .A3(new_n389), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n377), .A2(G200), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n401), .B2(KEYINPUT73), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT10), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT10), .B1(new_n377), .B2(G200), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT72), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n401), .A2(new_n410), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n392), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n313), .A2(new_n314), .ZN(new_n414));
  OAI21_X1  g0214(.A(G58), .B1(new_n219), .B2(new_n220), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n212), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(G20), .B1(G159), .B2(new_n301), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT7), .B1(new_n371), .B2(new_n216), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n251), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n250), .A2(new_n216), .A3(new_n251), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n420), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT78), .A3(G68), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n418), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n414), .B1(new_n430), .B2(KEYINPUT16), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT16), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n221), .B1(new_n427), .B2(new_n420), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT79), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n417), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g0235(.A(KEYINPUT79), .B(new_n221), .C1(new_n427), .C2(new_n420), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT80), .B(new_n432), .C1(new_n435), .C2(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n431), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n385), .B1(new_n263), .B2(G20), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n315), .B1(new_n385), .B2(new_n310), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G87), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n257), .A2(G1698), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G223), .B2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(new_n371), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n375), .B1(new_n447), .B2(new_n259), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT82), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n266), .B2(G232), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n265), .A2(KEYINPUT82), .A3(new_n337), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n448), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G190), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(G200), .B2(new_n452), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n443), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n441), .A2(KEYINPUT17), .A3(new_n443), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n441), .A2(new_n443), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n441), .A2(KEYINPUT81), .A3(new_n443), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n452), .A2(new_n347), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(G169), .B2(new_n452), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(KEYINPUT18), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT18), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n463), .A2(new_n470), .A3(new_n464), .A4(new_n467), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n366), .A2(new_n413), .A3(new_n469), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n263), .A2(G33), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n323), .B(new_n473), .C1(new_n297), .C2(new_n299), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT83), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n353), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n414), .A2(KEYINPUT83), .A3(new_n323), .A4(new_n473), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n252), .A2(new_n216), .A3(G68), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT19), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n216), .B1(new_n254), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G87), .B2(new_n206), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n304), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n300), .A2(new_n486), .B1(new_n310), .B2(new_n353), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n479), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT86), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n252), .A2(G244), .A3(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n490), .B(new_n491), .C1(new_n256), .C2(new_n222), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n259), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n269), .A2(G1), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n274), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n262), .C1(G250), .C2(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G179), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(G169), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n488), .A2(new_n489), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n498), .A2(G190), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(G200), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n476), .A2(G87), .A3(new_n478), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(new_n487), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n501), .A2(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n252), .A2(G257), .A3(G1698), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n252), .A2(G250), .A3(new_n255), .ZN(new_n510));
  INV_X1    g0310(.A(G294), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n249), .C2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n263), .B(G45), .C1(new_n268), .C2(KEYINPUT5), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .B1(KEYINPUT5), .B2(new_n268), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n494), .B(new_n515), .C1(KEYINPUT5), .C2(new_n268), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n259), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n259), .A2(new_n512), .B1(new_n517), .B2(G264), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n276), .A3(new_n516), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n310), .A2(new_n336), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT25), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n252), .A2(new_n216), .A3(G87), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT91), .B(KEYINPUT22), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n491), .B2(G20), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n216), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n336), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n526), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n414), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n526), .A2(new_n527), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n523), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n476), .A2(G107), .A3(new_n478), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n518), .A2(new_n519), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n521), .A2(new_n539), .A3(new_n540), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n336), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n484), .A2(new_n336), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n205), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(KEYINPUT6), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n428), .A2(G107), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n300), .B1(new_n484), .B2(new_n310), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n476), .A2(G97), .A3(new_n478), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(new_n255), .C1(new_n369), .C2(new_n370), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n252), .A2(KEYINPUT84), .A3(G250), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n262), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n517), .A2(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n519), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n344), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n565), .ZN(new_n569));
  INV_X1    g0369(.A(new_n567), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n347), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n553), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n565), .A2(new_n567), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n565), .B2(new_n567), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n552), .A4(new_n551), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n508), .A2(new_n543), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n474), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n315), .A2(KEYINPUT87), .A3(G116), .A4(new_n473), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n216), .A2(G116), .ZN(new_n583));
  AOI21_X1  g0383(.A(G20), .B1(new_n249), .B2(G97), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n558), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n311), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT88), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(KEYINPUT88), .A3(new_n587), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n309), .A2(G1), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n583), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n517), .A2(G270), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n252), .A2(G264), .A3(G1698), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n252), .A2(G257), .A3(new_n255), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n371), .A2(G303), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n259), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n600), .A3(new_n519), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n347), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n594), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT89), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT89), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n594), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(G200), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n595), .A2(new_n600), .A3(new_n519), .A4(G190), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(KEYINPUT90), .A3(new_n582), .A4(new_n593), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT90), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n594), .B2(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n601), .A2(G169), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n594), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n539), .A2(new_n540), .ZN(new_n622));
  AOI21_X1  g0422(.A(G169), .B1(new_n518), .B2(new_n519), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n347), .B2(new_n520), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n607), .A2(new_n615), .A3(new_n621), .A4(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n472), .A2(new_n577), .A3(new_n626), .ZN(G372));
  AND4_X1   g0427(.A1(new_n471), .A2(new_n366), .A3(new_n413), .A4(new_n469), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n488), .A2(new_n489), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n499), .A2(new_n500), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n502), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n553), .A2(new_n568), .A3(new_n571), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n507), .A2(new_n504), .A3(new_n503), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .ZN(new_n635));
  XNOR2_X1  g0435(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT94), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT94), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n635), .A2(new_n640), .A3(new_n631), .A4(new_n637), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n621), .A2(new_n607), .A3(new_n625), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n633), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n543), .A2(new_n576), .A3(new_n572), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n639), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n628), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT95), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT73), .ZN(new_n650));
  INV_X1    g0450(.A(new_n400), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n399), .B1(new_n388), .B2(new_n389), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n653), .B2(new_n397), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n654), .A2(new_n402), .A3(new_n404), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n655), .A2(KEYINPUT10), .B1(new_n409), .B2(new_n411), .ZN(new_n656));
  INV_X1    g0456(.A(new_n334), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n331), .B1(new_n657), .B2(new_n361), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n458), .A3(new_n459), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n466), .B1(new_n441), .B2(new_n443), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n660), .B(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n656), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n392), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n649), .A2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n605), .B1(new_n594), .B2(new_n602), .ZN(new_n668));
  INV_X1    g0468(.A(new_n606), .ZN(new_n669));
  INV_X1    g0469(.A(new_n620), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n619), .B1(new_n594), .B2(new_n616), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n592), .A2(new_n216), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(new_n594), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n594), .A2(new_n678), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n607), .A2(new_n621), .A3(new_n615), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n667), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n678), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n622), .A2(new_n624), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n622), .A2(new_n678), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n543), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(new_n625), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n678), .B1(new_n607), .B2(new_n621), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n625), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n209), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n213), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(new_n642), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n645), .A3(new_n615), .A4(new_n683), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n512), .A2(new_n259), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n517), .A2(G264), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n601), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n497), .A2(new_n347), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n573), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n705), .A2(new_n573), .A3(new_n706), .A4(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n541), .A2(new_n347), .A3(new_n497), .A4(new_n601), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n709), .B(new_n710), .C1(new_n573), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n678), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n667), .B1(new_n701), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n647), .A2(new_n683), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n642), .A2(new_n645), .B1(new_n502), .B2(new_n501), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n636), .B1(new_n508), .B2(new_n632), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n634), .A2(KEYINPUT26), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n678), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n718), .B1(new_n721), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n699), .B1(new_n728), .B2(G1), .ZN(G364));
  NAND3_X1  g0529(.A1(new_n679), .A2(new_n667), .A3(new_n681), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT97), .Z(new_n731));
  INV_X1    g0531(.A(new_n682), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n309), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n263), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n694), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n731), .A2(new_n732), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n679), .A2(new_n681), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G355), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n252), .A2(new_n209), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(G116), .B2(new_n209), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n246), .A2(G45), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n693), .A2(new_n252), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n269), .B2(new_n214), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT98), .ZN(new_n751));
  OAI21_X1  g0551(.A(G20), .B1(new_n751), .B2(G169), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n344), .A2(KEYINPUT98), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n275), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT99), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n741), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n736), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n216), .A2(KEYINPUT100), .A3(G190), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n347), .A2(G200), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT100), .B1(new_n216), .B2(G190), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G283), .A2(new_n766), .B1(new_n769), .B2(G329), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT102), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n216), .A2(new_n453), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n347), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G322), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n216), .A2(G190), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n773), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n763), .A2(new_n772), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n252), .B(new_n779), .C1(G303), .C2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n453), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n783), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(KEYINPUT33), .A2(G317), .ZN(new_n790));
  NAND2_X1  g0590(.A1(KEYINPUT33), .A2(G317), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n216), .B1(new_n767), .B2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n787), .B(new_n792), .C1(G294), .C2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n771), .A2(new_n782), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n793), .A2(new_n484), .ZN(new_n797));
  INV_X1    g0597(.A(new_n774), .ZN(new_n798));
  INV_X1    g0598(.A(new_n777), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G58), .A2(new_n798), .B1(new_n799), .B2(G77), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n320), .B2(new_n789), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n797), .B(new_n801), .C1(G50), .C2(new_n784), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n781), .A2(G87), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(KEYINPUT101), .A3(new_n252), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT101), .B1(new_n803), .B2(new_n252), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G107), .B2(new_n766), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n769), .A2(G159), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n796), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n761), .B1(new_n810), .B2(new_n758), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n742), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n738), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NAND2_X1  g0614(.A1(new_n360), .A2(new_n678), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n360), .A2(new_n349), .B1(new_n364), .B2(new_n815), .ZN(new_n816));
  AND4_X1   g0616(.A1(new_n360), .A2(new_n345), .A3(new_n348), .A4(new_n683), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT104), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n364), .A2(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n361), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT104), .ZN(new_n821));
  INV_X1    g0621(.A(new_n817), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n818), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n719), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n818), .A2(new_n823), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n683), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n647), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n626), .A2(new_n577), .A3(new_n678), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n715), .A2(new_n716), .ZN(new_n832));
  OAI21_X1  g0632(.A(G330), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT105), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n736), .B1(new_n830), .B2(new_n833), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n824), .A2(new_n739), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n758), .A2(new_n739), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n736), .B1(new_n840), .B2(G77), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n780), .A2(new_n336), .B1(new_n774), .B2(new_n511), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n252), .B(new_n842), .C1(G116), .C2(new_n799), .ZN(new_n843));
  INV_X1    g0643(.A(G303), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n785), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n797), .B(new_n845), .C1(G283), .C2(new_n788), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n769), .A2(G311), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n766), .A2(G87), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n252), .B1(new_n780), .B2(new_n387), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G58), .B2(new_n794), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n766), .A2(G68), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n768), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT103), .Z(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n798), .B1(new_n799), .B2(G159), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n784), .A2(G137), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n789), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT34), .Z(new_n860));
  OAI21_X1  g0660(.A(new_n849), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n841), .B1(new_n861), .B2(new_n758), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n837), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  XNOR2_X1  g0665(.A(new_n660), .B(new_n661), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n676), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  INV_X1    g0668(.A(new_n676), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n463), .A2(new_n464), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n456), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n468), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n441), .A2(new_n443), .A3(new_n455), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n431), .B1(KEYINPUT16), .B2(new_n430), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(new_n443), .B1(new_n466), .B2(new_n676), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n468), .A2(KEYINPUT18), .ZN(new_n879));
  INV_X1    g0679(.A(new_n460), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n471), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(new_n443), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n869), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n868), .B1(new_n874), .B2(new_n878), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n874), .A2(new_n878), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n331), .B(new_n334), .C1(new_n329), .C2(new_n683), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n330), .B(new_n678), .C1(new_n657), .C2(new_n292), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n638), .A2(KEYINPUT94), .B1(new_n645), .B2(new_n642), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n827), .B1(new_n893), .B2(new_n641), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n817), .B(KEYINPUT106), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(KEYINPUT107), .B(new_n867), .C1(new_n889), .C2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n456), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n441), .A2(KEYINPUT108), .A3(new_n443), .A4(new_n455), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n461), .A2(new_n467), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n870), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n874), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n460), .A2(KEYINPUT109), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT109), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n458), .A2(new_n908), .A3(new_n459), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n663), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n870), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n898), .B1(new_n913), .B2(new_n885), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n331), .A2(new_n678), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n883), .B1(new_n469), .B2(new_n471), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n874), .A2(new_n878), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n897), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n892), .ZN(new_n923));
  INV_X1    g0723(.A(new_n895), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n829), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n918), .A2(new_n919), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT107), .B1(new_n927), .B2(new_n867), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n721), .A2(new_n628), .A3(new_n727), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n665), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n929), .B(new_n931), .Z(new_n932));
  NAND2_X1  g0732(.A1(new_n701), .A2(new_n717), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n824), .B1(new_n890), .B2(new_n891), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n885), .B2(new_n888), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT40), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n908), .B1(new_n458), .B2(new_n459), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n866), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n870), .B1(new_n939), .B2(new_n909), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n441), .A2(KEYINPUT81), .A3(new_n443), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT81), .B1(new_n441), .B2(new_n443), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n872), .B1(new_n943), .B2(new_n467), .ZN(new_n944));
  AOI22_X1  g0744(.A1(KEYINPUT37), .A2(new_n904), .B1(new_n944), .B2(new_n870), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n868), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n919), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT40), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n936), .A2(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n628), .A3(new_n933), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n628), .A2(new_n933), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT40), .B1(new_n926), .B2(new_n935), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT40), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n946), .B2(new_n919), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(G330), .A3(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n932), .A2(new_n956), .B1(new_n263), .B2(new_n733), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT110), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n932), .A2(new_n956), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n963), .A2(G116), .A3(new_n217), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n214), .A2(G77), .A3(new_n415), .ZN(new_n967));
  INV_X1    g0767(.A(new_n201), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n320), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(G1), .A3(new_n309), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n962), .A2(new_n966), .A3(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n508), .B1(new_n507), .B2(new_n683), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n631), .A2(new_n507), .A3(new_n683), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n688), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT111), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n632), .A2(new_n678), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n553), .A2(new_n678), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n576), .A2(new_n572), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n982), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT111), .B1(new_n688), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n976), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(new_n976), .A3(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n981), .A2(new_n625), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n678), .B1(new_n990), .B2(new_n572), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n689), .A2(new_n687), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n982), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n994), .B2(KEYINPUT42), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(KEYINPUT42), .B2(new_n994), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n988), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n989), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n998), .A2(new_n999), .A3(new_n986), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n694), .B(KEYINPUT41), .Z(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT112), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n691), .A2(new_n1004), .A3(new_n982), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1004), .B1(new_n691), .B2(new_n982), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1007), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1009), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1010));
  OAI211_X1 g0810(.A(KEYINPUT44), .B(new_n984), .C1(new_n993), .C2(new_n684), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n691), .B2(new_n982), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1008), .A2(new_n1010), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n977), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1008), .A2(new_n1010), .A3(new_n688), .A4(new_n1014), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n689), .B(new_n687), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(new_n682), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n728), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n728), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1001), .B1(new_n1021), .B2(new_n735), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT113), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT113), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1001), .B(new_n1024), .C1(new_n1021), .C2(new_n735), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n972), .A2(new_n741), .A3(new_n973), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n238), .A2(new_n748), .B1(new_n209), .B2(new_n353), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n736), .B1(new_n760), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n793), .A2(new_n320), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G159), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n789), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G143), .B2(new_n784), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n780), .A2(new_n383), .B1(new_n777), .B2(new_n201), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n371), .B(new_n1035), .C1(G150), .C2(new_n798), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n766), .A2(G77), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n769), .A2(G137), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n780), .A2(new_n579), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1040), .A2(KEYINPUT46), .B1(new_n336), .B2(new_n793), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(KEYINPUT46), .B2(new_n1040), .ZN(new_n1042));
  INV_X1    g0842(.A(G283), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n371), .B1(new_n777), .B2(new_n1043), .C1(new_n789), .C2(new_n511), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G97), .B2(new_n766), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(KEYINPUT115), .B(G317), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n769), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1042), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n798), .A2(G303), .B1(G311), .B2(new_n784), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT114), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1039), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT47), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n758), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1029), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1027), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1026), .A2(new_n1057), .ZN(G387));
  NAND2_X1  g0858(.A1(new_n1019), .A2(new_n735), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n235), .A2(new_n269), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n351), .A2(G50), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT50), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n696), .B(new_n269), .C1(new_n320), .C2(new_n303), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n747), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1060), .B1(KEYINPUT116), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(KEYINPUT116), .B2(new_n1064), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(G107), .B2(new_n209), .C1(new_n696), .C2(new_n744), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n737), .B1(new_n1067), .B2(new_n759), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G97), .A2(new_n766), .B1(new_n769), .B2(G150), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n385), .B2(new_n789), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n780), .A2(new_n303), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n371), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n387), .B2(new_n774), .C1(new_n320), .C2(new_n777), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n794), .A2(new_n477), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n785), .B2(new_n1032), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n798), .A2(new_n1046), .B1(new_n799), .B2(G303), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n785), .B2(new_n775), .C1(new_n778), .C2(new_n789), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n780), .A2(new_n511), .B1(new_n793), .B2(new_n1043), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT117), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT49), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n371), .B1(new_n765), .B2(new_n579), .C1(new_n786), .C2(new_n768), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1085), .B2(KEYINPUT49), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1076), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n741), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1068), .B1(new_n1089), .B2(new_n1054), .C1(new_n687), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n728), .A2(new_n1019), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n694), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n728), .A2(new_n1019), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1059), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n1016), .A2(new_n735), .A3(new_n1017), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n785), .A2(new_n858), .B1(new_n774), .B2(new_n1032), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  OAI221_X1 g0898(.A(new_n252), .B1(new_n777), .B2(new_n351), .C1(new_n221), .C2(new_n780), .ZN(new_n1099));
  INV_X1    g0899(.A(G143), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n848), .B1(new_n1100), .B2(new_n768), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n789), .A2(new_n201), .B1(new_n303), .B2(new_n793), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n798), .A2(G311), .B1(G317), .B2(new_n784), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n371), .B1(new_n777), .B2(new_n511), .C1(new_n1043), .C2(new_n780), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n789), .A2(new_n844), .B1(new_n793), .B2(new_n579), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n336), .A2(new_n765), .B1(new_n768), .B2(new_n775), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT118), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n243), .A2(new_n748), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n759), .B1(new_n484), .B2(new_n209), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n736), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1110), .A2(new_n758), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n1111), .B2(new_n1114), .C1(new_n982), .C2(new_n1090), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1092), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1020), .A2(new_n694), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1096), .B(new_n1116), .C1(new_n1119), .C2(new_n1120), .ZN(G390));
  NAND4_X1  g0921(.A1(new_n933), .A2(G330), .A3(new_n826), .A4(new_n892), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n915), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n914), .A2(new_n920), .B1(new_n896), .B2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n678), .B(new_n824), .C1(new_n722), .C2(new_n725), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n892), .B1(new_n1126), .B2(new_n895), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n947), .A2(new_n1127), .A3(new_n1124), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1123), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n896), .A2(new_n1124), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n920), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT39), .B1(new_n946), .B2(new_n919), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n947), .A2(new_n1127), .A3(new_n1124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n1122), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n826), .C1(new_n831), .C2(new_n832), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n923), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n895), .B1(new_n726), .B2(new_n826), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1137), .A2(new_n1122), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1137), .A2(new_n1122), .B1(new_n829), .B2(new_n924), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n628), .A2(new_n718), .A3(KEYINPUT119), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n833), .B2(new_n472), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n930), .A2(new_n1145), .A3(new_n665), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1129), .A2(new_n1135), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n694), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(KEYINPUT120), .A3(new_n694), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1147), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1129), .A2(new_n1135), .A3(new_n735), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n739), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n737), .B1(new_n839), .B2(new_n385), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n789), .A2(new_n336), .B1(new_n303), .B2(new_n793), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G116), .A2(new_n798), .B1(new_n799), .B2(G97), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1161), .A2(new_n371), .A3(new_n803), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n852), .C1(new_n511), .C2(new_n768), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1160), .B(new_n1163), .C1(G283), .C2(new_n784), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT121), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n780), .A2(new_n858), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT53), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n1032), .B2(new_n793), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G137), .B2(new_n788), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n252), .B1(new_n774), .B2(new_n853), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n799), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1166), .A2(new_n1167), .B1(G128), .B2(new_n784), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G125), .A2(new_n769), .B1(new_n766), .B2(new_n968), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1169), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1165), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(KEYINPUT121), .B2(new_n1164), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1158), .B(new_n1159), .C1(new_n1054), .C2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1156), .A2(new_n1157), .A3(new_n1179), .ZN(G378));
  NOR2_X1   g0980(.A1(new_n391), .A2(new_n676), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n413), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n656), .B2(new_n392), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n949), .B2(G330), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n952), .A2(new_n954), .A3(new_n667), .A4(new_n1188), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1190), .A2(new_n1191), .B1(new_n928), .B2(new_n922), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n897), .A2(new_n921), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n948), .B1(new_n913), .B2(new_n885), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n933), .A2(new_n934), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n918), .B2(new_n919), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1194), .B(G330), .C1(new_n1196), .C2(KEYINPUT40), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1188), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n936), .A2(new_n937), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1199), .A2(G330), .A3(new_n1194), .A4(new_n1189), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n927), .A2(new_n867), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT107), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1193), .A2(new_n1198), .A3(new_n1200), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1192), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1146), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1148), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(KEYINPUT57), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT123), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT57), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1205), .A2(new_n1207), .A3(new_n1213), .A4(KEYINPUT57), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1209), .A2(new_n1212), .A3(new_n694), .A4(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1188), .A2(new_n739), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n784), .A2(G125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n789), .B2(new_n853), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n781), .A2(new_n1172), .B1(new_n799), .B2(G137), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n774), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(G150), .C2(new_n794), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n766), .A2(G159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1031), .B1(new_n785), .B2(new_n579), .C1(new_n484), .C2(new_n789), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n765), .A2(new_n383), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n371), .A2(new_n268), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n774), .A2(new_n336), .B1(new_n777), .B2(new_n353), .ZN(new_n1232));
  OR4_X1    g1032(.A1(new_n1071), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1229), .B(new_n1233), .C1(G283), .C2(new_n769), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT58), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1231), .B(new_n387), .C1(G33), .C2(G41), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1234), .A2(KEYINPUT58), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1228), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n758), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT122), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n839), .A2(new_n201), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1216), .A2(new_n736), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1205), .B2(new_n735), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1215), .A2(new_n1245), .ZN(G375));
  INV_X1    g1046(.A(new_n1002), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1154), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n734), .B(KEYINPUT124), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n736), .B1(new_n840), .B2(G68), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n780), .A2(new_n1032), .B1(new_n777), .B2(new_n858), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n371), .B(new_n1253), .C1(G137), .C2(new_n798), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1230), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n785), .A2(new_n853), .B1(new_n793), .B2(new_n387), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n788), .B2(new_n1172), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n769), .A2(G128), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1037), .A2(new_n371), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT125), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1074), .B1(new_n785), .B2(new_n511), .C1(new_n579), .C2(new_n789), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n780), .A2(new_n484), .B1(new_n777), .B2(new_n336), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G283), .B2(new_n798), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1263), .B(new_n1265), .C1(new_n844), .C2(new_n768), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1259), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1252), .B1(new_n1267), .B2(new_n758), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n892), .B2(new_n740), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1251), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1249), .A2(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G390), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n864), .ZN(new_n1274));
  OR4_X1    g1074(.A1(G396), .A2(new_n1274), .A3(G393), .A4(G381), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G387), .A2(new_n1275), .A3(G375), .A4(G378), .ZN(G407));
  AND3_X1   g1076(.A1(new_n1156), .A2(new_n1157), .A3(new_n1179), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n677), .A2(G213), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G407), .B(G213), .C1(G375), .C2(new_n1280), .ZN(G409));
  XNOR2_X1  g1081(.A(G393), .B(new_n813), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1023), .A2(new_n1025), .B1(new_n1027), .B2(new_n1056), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1273), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1285), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1289), .B(G390), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT61), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1215), .A2(G378), .A3(new_n1245), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1250), .B1(new_n1207), .B2(new_n1247), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1205), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1243), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1277), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1279), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1248), .B1(new_n1147), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1141), .A2(new_n1146), .A3(KEYINPUT60), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n694), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1271), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n864), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n864), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1279), .A2(G2897), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(G2897), .B(new_n1279), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1292), .B1(new_n1298), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1313), .B1(new_n1298), .B2(new_n1307), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1298), .A2(new_n1313), .A3(new_n1307), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1291), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1291), .B(new_n1292), .C1(new_n1298), .C2(new_n1311), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1298), .A2(new_n1307), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(KEYINPUT63), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1298), .A2(new_n1321), .A3(new_n1307), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1318), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT127), .B1(new_n1317), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1318), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1316), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1329), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1327), .B(new_n1328), .C1(new_n1330), .C2(new_n1291), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1324), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1277), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1293), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1307), .ZN(new_n1335));
  XOR2_X1   g1135(.A(new_n1335), .B(new_n1291), .Z(G402));
endmodule


