//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT64), .A2(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n194));
  AOI22_X1  g008(.A1(new_n191), .A2(new_n193), .B1(G128), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT64), .A2(G143), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(KEYINPUT65), .A3(G146), .A4(new_n198), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n189), .A2(new_n190), .A3(new_n188), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n192), .B2(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n199), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n195), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT11), .B1(new_n208), .B2(G137), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G137), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n208), .A2(KEYINPUT67), .A3(G137), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n208), .B2(G137), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n211), .A2(KEYINPUT68), .A3(G134), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n215), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G131), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT72), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n207), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n224), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT71), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n191), .A2(new_n193), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n189), .A2(new_n190), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n202), .B1(new_n238), .B2(G146), .ZN(new_n239));
  INV_X1    g053(.A(new_n199), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n233), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n203), .A2(new_n243), .A3(new_n233), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n237), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n213), .A2(new_n217), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n219), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n230), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n202), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n197), .A2(new_n198), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(new_n188), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT66), .B(new_n232), .C1(new_n252), .C2(new_n199), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n243), .B1(new_n203), .B2(new_n233), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n248), .B(new_n236), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n229), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n258));
  INV_X1    g072(.A(G119), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G119), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n262), .A3(G116), .ZN(new_n263));
  INV_X1    g077(.A(G116), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G119), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT2), .B(G113), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n266), .B2(new_n267), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n267), .ZN(new_n273));
  INV_X1    g087(.A(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT73), .A3(new_n269), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n257), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n277), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n229), .C1(new_n249), .C2(new_n256), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(KEYINPUT78), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n228), .A2(new_n227), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n282), .A2(new_n207), .A3(new_n225), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n255), .A2(KEYINPUT71), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n242), .A2(new_n244), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n285), .A2(new_n230), .A3(new_n248), .A4(new_n236), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  OR3_X1    g101(.A1(new_n287), .A2(KEYINPUT78), .A3(new_n279), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n281), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT74), .B(KEYINPUT27), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT75), .ZN(new_n291));
  INV_X1    g105(.A(G237), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(G210), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n291), .B(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G101), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n229), .A2(new_n255), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n229), .A2(new_n301), .A3(new_n255), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n279), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n289), .A2(KEYINPUT29), .A3(new_n298), .A4(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n207), .A2(new_n228), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n255), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n275), .A2(new_n269), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n280), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g127(.A(KEYINPUT76), .B(new_n304), .C1(new_n280), .C2(new_n310), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n313), .A2(new_n297), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n283), .B(new_n277), .C1(new_n284), .C2(new_n286), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n308), .A2(KEYINPUT30), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n287), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(new_n309), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n316), .B1(new_n322), .B2(new_n298), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n187), .B(new_n306), .C1(new_n315), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT32), .ZN(new_n326));
  NOR2_X1   g140(.A1(G472), .A2(G902), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n318), .B1(new_n257), .B2(KEYINPUT30), .ZN(new_n328));
  INV_X1    g142(.A(new_n309), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n298), .B(new_n280), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT31), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT31), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n322), .A2(new_n332), .A3(new_n298), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n277), .B1(new_n299), .B2(KEYINPUT77), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT28), .B1(new_n335), .B2(new_n302), .ZN(new_n336));
  INV_X1    g150(.A(new_n310), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT28), .B1(new_n317), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n311), .A2(new_n312), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n298), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n326), .B(new_n327), .C1(new_n334), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n297), .B1(new_n313), .B2(new_n314), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n331), .A3(new_n333), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n326), .B1(new_n345), .B2(new_n327), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n325), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n350), .A2(KEYINPUT16), .A3(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(G146), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G146), .B1(new_n349), .B2(new_n351), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n260), .A2(new_n262), .A3(G128), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n259), .B2(G128), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT24), .B(G110), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n260), .A2(new_n262), .ZN(new_n362));
  INV_X1    g176(.A(G128), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT79), .B1(new_n356), .B2(KEYINPUT23), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(KEYINPUT23), .A3(G119), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G110), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n360), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT80), .B(G110), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n368), .B(new_n372), .C1(new_n365), .C2(new_n366), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n357), .A2(new_n358), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT81), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n188), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT82), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(new_n352), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT81), .B1(new_n373), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT22), .B(G137), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n293), .A2(G221), .A3(G234), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT83), .Z(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n371), .B(new_n384), .C1(new_n379), .C2(new_n380), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n187), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n386), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n387), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(KEYINPUT84), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(G234), .B2(new_n187), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n395), .A3(new_n389), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n394), .A2(G902), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n387), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n377), .B1(new_n188), .B2(new_n348), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n292), .A2(new_n293), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G143), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n251), .B2(new_n405), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT91), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  OAI22_X1  g223(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n214), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n251), .A2(new_n405), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n214), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(KEYINPUT91), .A3(new_n412), .A4(new_n406), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(G131), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n214), .A3(new_n406), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n348), .B(KEYINPUT19), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n188), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n352), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  INV_X1    g237(.A(G104), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n407), .A2(KEYINPUT17), .A3(G131), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n355), .B(new_n428), .C1(new_n418), .C2(KEYINPUT17), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n415), .A3(new_n425), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT20), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n435), .A3(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(new_n430), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n425), .B1(new_n429), .B2(new_n415), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n187), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT92), .B(G475), .Z(new_n440));
  AOI22_X1  g254(.A1(new_n434), .A2(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n197), .A2(G128), .A3(new_n198), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n363), .A2(G143), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n208), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(G107), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AND4_X1   g261(.A1(KEYINPUT93), .A2(new_n442), .A3(KEYINPUT13), .A4(new_n443), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n449));
  OAI21_X1  g263(.A(G134), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n444), .B(new_n447), .C1(new_n448), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n446), .B1(new_n453), .B2(KEYINPUT14), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(G116), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n264), .A2(G122), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n454), .A2(KEYINPUT94), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT94), .B1(new_n454), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n445), .A2(new_n446), .ZN(new_n462));
  INV_X1    g276(.A(new_n444), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n208), .B1(new_n442), .B2(new_n443), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n451), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT9), .B(G234), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n467), .A2(new_n393), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n451), .B(new_n468), .C1(new_n461), .C2(new_n465), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(KEYINPUT95), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n473), .A3(new_n469), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n187), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n475), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(G952), .A3(new_n293), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n441), .A2(new_n479), .A3(KEYINPUT96), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT96), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n439), .A2(new_n440), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n491));
  INV_X1    g305(.A(new_n432), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT20), .B(new_n492), .C1(new_n427), .C2(new_n430), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n490), .B(new_n487), .C1(new_n491), .C2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n489), .B1(new_n494), .B2(new_n478), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G210), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n501));
  XNOR2_X1  g315(.A(G110), .B(G122), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n446), .A2(G104), .ZN(new_n505));
  AND2_X1   g319(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT87), .B(G101), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n424), .A2(G107), .ZN(new_n509));
  NOR2_X1   g323(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(G104), .A3(new_n446), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G101), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(KEYINPUT4), .A3(G101), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n516), .A2(new_n517), .B1(new_n269), .B2(new_n275), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n274), .A2(new_n263), .A3(new_n265), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n263), .A2(KEYINPUT5), .A3(new_n265), .ZN(new_n520));
  OAI21_X1  g334(.A(G113), .B1(new_n263), .B2(KEYINPUT5), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n505), .A2(new_n509), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G101), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n501), .B(new_n503), .C1(new_n518), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT90), .ZN(new_n528));
  AOI22_X1  g342(.A1(KEYINPUT4), .A2(new_n512), .B1(new_n514), .B2(G101), .ZN(new_n529));
  INV_X1    g343(.A(new_n517), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n309), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n526), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n501), .A4(new_n503), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n207), .A2(new_n350), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n245), .B2(new_n350), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(G224), .A3(new_n293), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n236), .B1(new_n253), .B2(new_n254), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G125), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n293), .A2(G224), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n503), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n516), .A2(new_n517), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n526), .B1(new_n546), .B2(new_n309), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n502), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT6), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n536), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n522), .B(new_n525), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n502), .B(KEYINPUT8), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n547), .A2(new_n502), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n541), .A2(KEYINPUT7), .A3(new_n542), .A4(new_n537), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n538), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n539), .A2(new_n553), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n187), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n500), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n536), .A2(new_n544), .A3(new_n549), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n560), .A2(new_n187), .A3(new_n499), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n498), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G221), .B1(new_n467), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G469), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n293), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n512), .A2(new_n524), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT10), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n363), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n203), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n205), .B1(new_n252), .B2(new_n199), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n570), .B(new_n571), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT10), .B1(new_n207), .B2(new_n525), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n245), .A2(new_n546), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n248), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT88), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n546), .A2(new_n285), .A3(new_n236), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n248), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n581), .A3(new_n578), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n569), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT89), .A3(new_n569), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n570), .A2(new_n195), .A3(new_n574), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n204), .B1(new_n251), .B2(new_n188), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n252), .B(new_n199), .C1(new_n590), .C2(new_n363), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n203), .A2(new_n206), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n525), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n248), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT12), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n207), .A2(new_n525), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n578), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT12), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n588), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT89), .B1(new_n586), .B2(new_n569), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n565), .B(new_n187), .C1(new_n587), .C2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n568), .B1(new_n577), .B2(new_n578), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n599), .A2(KEYINPUT12), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n595), .B(new_n578), .C1(new_n597), .C2(new_n598), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n586), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n585), .A2(new_n606), .B1(new_n568), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G469), .B1(new_n610), .B2(G902), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n564), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n496), .A2(new_n562), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n347), .A2(new_n403), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(new_n508), .Z(G3));
  NAND2_X1  g429(.A1(new_n605), .A2(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n563), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n401), .A2(new_n402), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G472), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n345), .B2(new_n187), .ZN(new_n620));
  INV_X1    g434(.A(new_n327), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n331), .A2(new_n333), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n344), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n562), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n472), .A2(new_n627), .A3(new_n474), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n470), .A2(KEYINPUT33), .A3(new_n471), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n476), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n475), .A2(KEYINPUT97), .A3(new_n476), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT97), .B1(new_n475), .B2(new_n476), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n490), .B1(new_n491), .B2(new_n493), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n626), .A2(new_n486), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n625), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NOR2_X1   g455(.A1(new_n479), .A2(new_n636), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n562), .A2(new_n487), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n385), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n381), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n399), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n397), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n396), .A2(new_n394), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n653), .A2(new_n392), .B1(new_n399), .B2(new_n648), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n613), .A3(new_n624), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  XNOR2_X1  g474(.A(new_n481), .B(KEYINPUT99), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n662), .B1(new_n663), .B2(new_n484), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n617), .A2(new_n626), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n347), .A2(new_n657), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n664), .B(KEYINPUT39), .Z(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n612), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n559), .A2(new_n561), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n559), .A2(KEYINPUT38), .A3(new_n561), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n636), .A2(new_n478), .A3(new_n497), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n672), .A2(new_n677), .A3(new_n650), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n281), .A2(new_n297), .A3(new_n288), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n330), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT100), .ZN(new_n682));
  AOI21_X1  g496(.A(G902), .B1(new_n681), .B2(KEYINPUT100), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI22_X1  g498(.A1(new_n684), .A2(new_n619), .B1(new_n343), .B2(new_n346), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n612), .A2(new_n671), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n670), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n251), .ZN(G45));
  NOR2_X1   g503(.A1(new_n637), .A2(new_n664), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n691), .A2(new_n617), .A3(new_n626), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n347), .A2(new_n657), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  INV_X1    g508(.A(new_n402), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n327), .B1(new_n334), .B2(new_n341), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT32), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n342), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n697), .B1(new_n700), .B2(new_n325), .ZN(new_n701));
  INV_X1    g515(.A(new_n605), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n579), .A2(new_n584), .B1(new_n578), .B2(new_n577), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n703), .A2(new_n569), .B1(new_n602), .B2(new_n603), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n565), .B1(new_n704), .B2(new_n187), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n702), .A2(new_n705), .A3(new_n564), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n638), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  AND2_X1   g524(.A1(new_n643), .A2(new_n706), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  NAND3_X1  g527(.A1(new_n706), .A2(KEYINPUT101), .A3(new_n562), .ZN(new_n714));
  INV_X1    g528(.A(new_n705), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n562), .A3(new_n563), .A4(new_n605), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n347), .A3(new_n496), .A4(new_n657), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AOI21_X1  g535(.A(new_n298), .B1(new_n289), .B2(new_n305), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n327), .B1(new_n334), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n187), .B1(new_n334), .B2(new_n341), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G472), .ZN(new_n727));
  OAI211_X1 g541(.A(KEYINPUT102), .B(new_n327), .C1(new_n334), .C2(new_n722), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n397), .A2(new_n400), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n678), .B1(new_n559), .B2(new_n561), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n706), .A2(new_n487), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND4_X1  g549(.A1(new_n729), .A2(new_n719), .A3(new_n650), .A4(new_n690), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  AOI22_X1  g551(.A1(new_n699), .A2(new_n342), .B1(G472), .B2(new_n324), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT104), .B1(new_n673), .B2(new_n498), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n559), .A2(new_n740), .A3(new_n497), .A4(new_n561), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT103), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n610), .B2(G469), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n564), .B1(new_n605), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n739), .A2(new_n690), .A3(new_n741), .A4(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n738), .A2(new_n730), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n739), .A2(new_n741), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n347), .A2(new_n403), .A3(new_n751), .A4(new_n746), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n690), .A2(new_n749), .ZN(new_n753));
  OAI22_X1  g567(.A1(new_n748), .A2(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n214), .ZN(G33));
  INV_X1    g569(.A(new_n666), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n701), .A2(new_n756), .A3(new_n751), .A4(new_n746), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  AND3_X1   g572(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n475), .A2(new_n476), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n759), .B1(new_n762), .B2(new_n632), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n763), .B2(new_n636), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n635), .A2(new_n441), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n654), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n620), .B2(new_n623), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n750), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n768), .B(KEYINPUT44), .C1(new_n620), .C2(new_n623), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n586), .A2(new_n569), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n579), .B2(new_n584), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n569), .B1(new_n601), .B2(new_n586), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n583), .B1(new_n582), .B2(new_n248), .ZN(new_n778));
  AOI211_X1 g592(.A(KEYINPUT88), .B(new_n578), .C1(new_n580), .C2(new_n581), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n606), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n609), .A2(new_n568), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT45), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(new_n782), .A3(G469), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n743), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n702), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n564), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT105), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n788), .A2(new_n789), .A3(new_n671), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n789), .B1(new_n788), .B2(new_n671), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n771), .B(new_n772), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NOR3_X1   g607(.A1(new_n403), .A2(new_n691), .A3(new_n750), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n796), .B(new_n564), .C1(new_n786), .C2(new_n787), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n794), .B(new_n738), .C1(new_n795), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NAND2_X1  g613(.A1(new_n715), .A2(new_n605), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT49), .Z(new_n801));
  AOI21_X1  g615(.A(new_n619), .B1(new_n682), .B2(new_n683), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n699), .B2(new_n342), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n763), .A2(new_n636), .A3(new_n498), .A4(new_n564), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n677), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n801), .A2(new_n731), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n725), .A2(new_n727), .A3(new_n731), .A4(new_n728), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n767), .A2(new_n661), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n751), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n800), .A2(new_n563), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n795), .A2(new_n797), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT108), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n816));
  INV_X1    g630(.A(new_n797), .ZN(new_n817));
  INV_X1    g631(.A(new_n813), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n751), .A4(new_n811), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n715), .A2(new_n563), .A3(new_n605), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT114), .B1(new_n750), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n706), .A2(new_n825), .A3(new_n741), .A4(new_n739), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n697), .A2(new_n481), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n763), .A2(new_n441), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n827), .A2(new_n803), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT115), .B1(new_n827), .B2(new_n809), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n835), .B(new_n810), .C1(new_n824), .C2(new_n826), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n650), .B(new_n729), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n832), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n822), .A2(new_n833), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT109), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n559), .A2(KEYINPUT38), .A3(new_n561), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT38), .B1(new_n559), .B2(new_n561), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n498), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n843), .B2(new_n823), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n677), .A2(new_n706), .A3(KEYINPUT109), .A4(new_n498), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n811), .A2(new_n846), .A3(KEYINPUT50), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n811), .A2(new_n846), .A3(KEYINPUT110), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n724), .A2(new_n723), .B1(new_n726), .B2(G472), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n731), .A3(new_n728), .A4(new_n809), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n845), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n855));
  AOI21_X1  g669(.A(KEYINPUT112), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  INV_X1    g671(.A(new_n855), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n857), .B(new_n858), .C1(new_n848), .C2(new_n853), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n847), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n839), .B1(new_n860), .B2(KEYINPUT113), .ZN(new_n861));
  INV_X1    g675(.A(new_n847), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT110), .B1(new_n811), .B2(new_n846), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n851), .A2(new_n852), .A3(new_n849), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n855), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n857), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n837), .A2(new_n833), .A3(new_n838), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT51), .B1(new_n812), .B2(new_n814), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n860), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n827), .A2(new_n803), .A3(new_n828), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(new_n637), .ZN(new_n877));
  INV_X1    g691(.A(G952), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n878), .B(G953), .C1(new_n811), .C2(new_n719), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT117), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n730), .B1(new_n700), .B2(new_n325), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n834), .B2(new_n836), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n879), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n875), .A2(new_n880), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n807), .B1(new_n871), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(new_n822), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n872), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n868), .B2(new_n869), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n860), .A2(KEYINPUT113), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n875), .A2(new_n887), .A3(new_n880), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT118), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n347), .B(new_n403), .C1(new_n707), .C2(new_n711), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n720), .A3(new_n734), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n618), .B(new_n624), .C1(new_n638), .C2(new_n643), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n614), .A2(new_n902), .A3(new_n658), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n614), .A2(new_n902), .A3(new_n658), .A4(KEYINPUT106), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n739), .A2(new_n741), .A3(new_n746), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n729), .A2(new_n650), .A3(new_n690), .A4(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n636), .A2(new_n478), .A3(new_n664), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n739), .A2(new_n741), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT107), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n617), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n739), .A2(KEYINPUT107), .A3(new_n741), .A4(new_n910), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n347), .A3(new_n657), .A4(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n909), .B(new_n915), .C1(new_n666), .C2(new_n752), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(new_n754), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n654), .A2(new_n732), .A3(new_n665), .A4(new_n746), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n685), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n736), .A2(new_n668), .A3(new_n693), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT52), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n725), .A2(new_n727), .A3(new_n650), .A4(new_n728), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n691), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n656), .B1(new_n700), .B2(new_n325), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n923), .A2(new_n719), .B1(new_n924), .B2(new_n667), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT52), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n693), .A4(new_n919), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n907), .A2(new_n917), .A3(new_n921), .A4(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n920), .A2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n899), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n921), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(KEYINPUT53), .A3(new_n907), .A4(new_n917), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n898), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT53), .B1(new_n928), .B2(new_n929), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n899), .A3(new_n907), .A4(new_n917), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT54), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n889), .A2(new_n897), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(G952), .A2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n806), .B1(new_n939), .B2(new_n940), .ZN(G75));
  NAND4_X1  g755(.A1(new_n935), .A2(G210), .A3(G902), .A4(new_n936), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n536), .A2(new_n549), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n544), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT55), .Z(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(KEYINPUT56), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n942), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n942), .B2(new_n948), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n293), .A2(G952), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(G51));
  NAND2_X1  g766(.A1(new_n935), .A2(new_n936), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n898), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n954), .A2(new_n937), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n743), .B(KEYINPUT57), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n704), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n953), .A2(new_n187), .A3(new_n783), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n951), .B1(new_n957), .B2(new_n958), .ZN(G54));
  NOR2_X1   g773(.A1(new_n953), .A2(new_n187), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  INV_X1    g775(.A(new_n431), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n951), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(KEYINPUT58), .A3(G475), .A4(new_n431), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G60));
  AND2_X1   g779(.A1(new_n628), .A2(new_n629), .ZN(new_n966));
  NAND2_X1  g780(.A1(G478), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT59), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n955), .A2(new_n969), .B1(G952), .B2(new_n293), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n934), .A2(new_n937), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n971), .B2(new_n968), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT60), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n935), .A2(new_n936), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n386), .A2(new_n387), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n951), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n935), .A2(new_n648), .A3(new_n936), .A4(new_n975), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(KEYINPUT120), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(KEYINPUT120), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(KEYINPUT61), .B(new_n978), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  INV_X1    g800(.A(G224), .ZN(new_n987));
  OAI21_X1  g801(.A(G953), .B1(new_n485), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT121), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n907), .B(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n990), .B2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n943), .B1(G898), .B2(new_n293), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n347), .A2(new_n731), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT42), .B1(new_n994), .B2(new_n747), .ZN(new_n995));
  INV_X1    g809(.A(new_n753), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n701), .A2(new_n751), .A3(new_n746), .A4(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n995), .A2(new_n997), .A3(new_n757), .A4(new_n798), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n736), .A2(new_n668), .A3(new_n693), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n771), .A2(new_n772), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n881), .A2(new_n732), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n790), .A2(new_n791), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1000), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n999), .A2(new_n1006), .A3(KEYINPUT124), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n771), .A2(new_n772), .B1(new_n881), .B2(new_n732), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n693), .B(new_n925), .C1(new_n1009), .C2(new_n1004), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1008), .B1(new_n1010), .B2(new_n998), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n1011), .A3(new_n293), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n328), .B(new_n419), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(G900), .B2(G953), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n637), .B1(new_n479), .B2(new_n636), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT122), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n701), .A2(new_n686), .A3(new_n751), .A4(new_n1016), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n792), .A2(new_n798), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n925), .A2(new_n1019), .A3(new_n688), .A4(new_n693), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n736), .A2(new_n688), .A3(new_n668), .A4(new_n693), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1018), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n293), .ZN(new_n1025));
  AOI22_X1  g839(.A1(new_n1012), .A2(new_n1014), .B1(new_n1025), .B2(new_n1013), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT123), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1026), .B(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  NOR2_X1   g846(.A1(new_n907), .A2(new_n989), .ZN(new_n1033));
  AOI211_X1 g847(.A(KEYINPUT121), .B(new_n901), .C1(new_n905), .C2(new_n906), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n322), .A2(new_n297), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n951), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1032), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n322), .A2(new_n297), .ZN(new_n1042));
  AOI21_X1  g856(.A(KEYINPUT125), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT125), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1042), .ZN(new_n1045));
  AOI211_X1 g859(.A(new_n1044), .B(new_n1045), .C1(new_n1040), .C2(new_n1032), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1039), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g861(.A(KEYINPUT126), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n930), .A2(new_n933), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1032), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1038), .A2(new_n1042), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1048), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1051), .ZN(new_n1053));
  AOI211_X1 g867(.A(KEYINPUT126), .B(new_n1053), .C1(new_n930), .C2(new_n933), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(KEYINPUT127), .B1(new_n1047), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n905), .A2(new_n906), .ZN(new_n1057));
  INV_X1    g871(.A(new_n901), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n917), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1059), .A2(new_n899), .A3(new_n931), .ZN(new_n1060));
  INV_X1    g874(.A(new_n929), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n932), .A2(new_n907), .A3(new_n917), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1060), .B1(new_n899), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g877(.A(KEYINPUT126), .B1(new_n1063), .B2(new_n1053), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1049), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(KEYINPUT127), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1050), .B1(new_n990), .B2(new_n1023), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1044), .B1(new_n1068), .B2(new_n1045), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1041), .A2(KEYINPUT125), .A3(new_n1042), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g885(.A1(new_n1066), .A2(new_n1067), .A3(new_n1071), .A4(new_n1039), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1056), .A2(new_n1072), .ZN(G57));
endmodule


