//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n209), .B1(new_n211), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G68), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n226), .B1(G238), .B2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT67), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n231), .B(new_n232), .C1(new_n228), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n206), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n220), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n235), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G222), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G223), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n261), .B(new_n262), .C1(G77), .C2(new_n257), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n265), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(G226), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G179), .ZN(new_n271));
  XOR2_X1   g0071(.A(new_n271), .B(KEYINPUT70), .Z(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT8), .A2(G58), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT68), .B(G58), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(KEYINPUT8), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n204), .A3(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n222), .A2(new_n212), .A3(new_n213), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n277), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n210), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n280), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n203), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  MUX2_X1   g0090(.A(new_n287), .B(new_n290), .S(G50), .Z(new_n291));
  NAND3_X1  g0091(.A1(new_n284), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n270), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n272), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n227), .A2(new_n204), .ZN(new_n297));
  INV_X1    g0097(.A(new_n278), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n204), .A2(G33), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n298), .A2(new_n222), .B1(new_n299), .B2(new_n224), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n282), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT11), .ZN(new_n302));
  INV_X1    g0102(.A(new_n287), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT73), .B1(new_n303), .B2(new_n282), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n287), .A2(new_n305), .A3(new_n210), .A4(new_n281), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n304), .A2(G68), .A3(new_n289), .A4(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(KEYINPUT12), .A2(G68), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n287), .A2(new_n308), .A3(KEYINPUT77), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT12), .B1(new_n227), .B2(new_n287), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT77), .B1(new_n287), .B2(new_n308), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n307), .A2(new_n312), .A3(KEYINPUT78), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n302), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n223), .A2(new_n259), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n259), .A2(G232), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n257), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n262), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n266), .B1(G238), .B2(new_n268), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n262), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n320), .B2(new_n321), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n262), .A2(new_n264), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n267), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(G238), .A3(new_n265), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT13), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT14), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(G169), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n326), .A2(new_n333), .A3(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n335), .B1(new_n334), .B2(G169), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n317), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n296), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g0142(.A(KEYINPUT8), .B(G58), .Z(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n344), .A2(new_n345), .B1(new_n299), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n282), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n303), .A2(new_n224), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G232), .A2(G1698), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n259), .A2(G238), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n257), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G107), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G107), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n354), .B(new_n262), .C1(new_n257), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n266), .B1(G244), .B2(new_n268), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n304), .A2(G77), .A3(new_n289), .A4(new_n306), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT74), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(G190), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n351), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(G169), .B1(new_n360), .B2(new_n361), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n362), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n349), .A3(new_n350), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT75), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n292), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n270), .A2(G200), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n284), .A2(KEYINPUT9), .A3(new_n286), .A4(new_n291), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n263), .A2(new_n269), .A3(G190), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n378), .B2(KEYINPUT76), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n381), .B(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n324), .B1(new_n323), .B2(new_n325), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n328), .A2(new_n332), .A3(KEYINPUT13), .ZN(new_n387));
  OAI21_X1  g0187(.A(G200), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n326), .A2(new_n333), .A3(G190), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n390), .B2(new_n317), .ZN(new_n391));
  INV_X1    g0191(.A(new_n317), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n392), .A2(new_n388), .A3(KEYINPUT79), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n342), .A2(new_n375), .A3(new_n384), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n253), .A2(KEYINPUT80), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n399), .A3(G33), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n256), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI211_X1 g0203(.A(KEYINPUT7), .B(G20), .C1(new_n400), .C2(new_n256), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n256), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(G33), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT7), .B1(new_n408), .B2(G20), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n401), .A2(new_n402), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT81), .A4(G68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT82), .ZN(new_n413));
  NOR2_X1   g0213(.A1(KEYINPUT66), .A2(G68), .ZN(new_n414));
  AND2_X1   g0214(.A1(KEYINPUT66), .A2(G68), .ZN(new_n415));
  AND2_X1   g0215(.A1(KEYINPUT68), .A2(G58), .ZN(new_n416));
  NOR2_X1   g0216(.A1(KEYINPUT68), .A2(G58), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n414), .A2(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n204), .B1(new_n418), .B2(new_n214), .ZN(new_n419));
  INV_X1    g0219(.A(G159), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n298), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n413), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n227), .A2(new_n274), .B1(new_n212), .B2(new_n213), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT82), .B(new_n423), .C1(new_n424), .C2(new_n204), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n422), .A2(KEYINPUT16), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n412), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n428));
  INV_X1    g0228(.A(new_n227), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT84), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n402), .C1(new_n257), .C2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(G20), .B1(new_n254), .B2(new_n256), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT84), .B1(new_n432), .B2(KEYINPUT7), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(KEYINPUT85), .B(new_n254), .C1(new_n407), .C2(G33), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n397), .A2(new_n399), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT85), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n255), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n429), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n422), .A2(new_n425), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n428), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n427), .A2(new_n442), .A3(new_n282), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n275), .A2(new_n303), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n275), .B2(new_n290), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n266), .B1(G232), .B2(new_n268), .ZN(new_n447));
  NOR2_X1   g0247(.A1(G223), .A2(G1698), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n448), .B1(new_n223), .B2(G1698), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n408), .A2(new_n449), .B1(G33), .B2(G87), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n447), .B1(new_n327), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n363), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G190), .B2(new_n451), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n443), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n288), .B1(new_n412), .B2(new_n426), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n445), .B1(new_n457), .B2(new_n442), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(KEYINPUT17), .A3(new_n453), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n443), .A2(new_n446), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n408), .A2(new_n449), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G87), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n327), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n268), .A2(G232), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n330), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n293), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT86), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n447), .B(new_n370), .C1(new_n327), .C2(new_n450), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(new_n472), .A3(KEYINPUT18), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT18), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n470), .A2(new_n471), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n458), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT87), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(KEYINPUT87), .B(new_n474), .C1(new_n458), .C2(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n460), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n395), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT22), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n400), .A2(new_n204), .A3(G87), .A4(new_n256), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT95), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n408), .A2(KEYINPUT95), .A3(new_n204), .A4(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n254), .A2(new_n256), .ZN(new_n490));
  INV_X1    g0290(.A(G87), .ZN(new_n491));
  NOR4_X1   g0291(.A1(new_n490), .A2(KEYINPUT22), .A3(G20), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n495));
  INV_X1    g0295(.A(new_n359), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n495), .B1(new_n497), .B2(KEYINPUT23), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT89), .B(G116), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G33), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT96), .B1(new_n501), .B2(G20), .ZN(new_n502));
  OR4_X1    g0302(.A1(KEYINPUT96), .A2(new_n499), .A3(G20), .A4(new_n255), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n483), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n492), .B1(new_n487), .B2(new_n488), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT24), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n282), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n203), .A2(G33), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n288), .A2(new_n287), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT25), .B1(new_n303), .B2(new_n355), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n355), .ZN(new_n515));
  AOI22_X1  g0315(.A1(G107), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G250), .A2(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(G257), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(G1698), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n408), .A2(new_n520), .B1(G33), .B2(G294), .ZN(new_n521));
  INV_X1    g0321(.A(G264), .ZN(new_n522));
  XNOR2_X1  g0322(.A(KEYINPUT5), .B(G41), .ZN(new_n523));
  INV_X1    g0323(.A(G45), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G1), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n327), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n521), .A2(new_n327), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n526), .A2(new_n264), .A3(new_n262), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n528), .A2(G179), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n532), .B2(new_n293), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n517), .A2(KEYINPUT97), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n494), .A2(new_n504), .A3(new_n483), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT24), .B1(new_n506), .B2(new_n507), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n288), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n516), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n531), .A2(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n532), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n509), .A2(new_n542), .A3(new_n516), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n400), .A2(new_n256), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n259), .A2(G244), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n548), .A2(new_n546), .B1(new_n550), .B2(new_n259), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n257), .A2(new_n551), .B1(G33), .B2(G283), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n327), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n329), .A2(new_n525), .A3(new_n523), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n519), .B2(new_n527), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n553), .A2(new_n555), .A3(G179), .ZN(new_n556));
  INV_X1    g0356(.A(new_n527), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n529), .B1(G257), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n549), .A2(new_n552), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n327), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n556), .B1(new_n293), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n496), .B1(new_n434), .B2(new_n439), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G97), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n564), .A2(new_n566), .A3(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n568), .A2(new_n204), .B1(new_n224), .B2(new_n298), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n282), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n303), .A2(new_n566), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n511), .B2(new_n566), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n561), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n553), .A2(new_n555), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT88), .B1(new_n576), .B2(G190), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT88), .ZN(new_n578));
  INV_X1    g0378(.A(G190), .ZN(new_n579));
  NOR4_X1   g0379(.A1(new_n553), .A2(new_n555), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n553), .B2(new_n555), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n570), .A2(new_n573), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n575), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT94), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G257), .A2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n522), .B2(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n408), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n490), .A2(G303), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n327), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G270), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n554), .B1(new_n591), .B2(new_n527), .ZN(new_n592));
  OAI21_X1  g0392(.A(G169), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n304), .A2(G116), .A3(new_n306), .A4(new_n510), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n499), .A2(new_n303), .ZN(new_n595));
  AOI21_X1  g0395(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G283), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n210), .B2(new_n281), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n499), .A2(G20), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT20), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT20), .B1(new_n598), .B2(new_n599), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n594), .B(new_n595), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n585), .B1(new_n593), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n590), .A2(new_n592), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n603), .C1(new_n363), .C2(new_n606), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n590), .A2(new_n592), .A3(new_n370), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n602), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n585), .B(new_n611), .C1(new_n593), .C2(new_n603), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n605), .A2(new_n608), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n584), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n525), .A2(new_n264), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n550), .B1(new_n524), .B2(G1), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n327), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(G238), .A2(G1698), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n225), .B2(G1698), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n408), .A2(new_n619), .B1(G33), .B2(new_n500), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n327), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n293), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n370), .B(new_n617), .C1(new_n620), .C2(new_n327), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n400), .A2(new_n204), .A3(G68), .A4(new_n256), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT19), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n356), .A2(new_n358), .A3(new_n491), .A4(new_n566), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n321), .A2(new_n204), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n299), .A2(KEYINPUT19), .A3(new_n566), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n282), .B1(new_n303), .B2(new_n346), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT91), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n346), .B(KEYINPUT90), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n511), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT90), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n346), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n512), .A3(KEYINPUT91), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT92), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n632), .A2(new_n639), .A3(KEYINPUT92), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n624), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n617), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n408), .A2(new_n619), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n501), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n262), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G190), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n512), .A2(G87), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n621), .A2(G200), .ZN(new_n651));
  AND4_X1   g0451(.A1(new_n632), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT93), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n624), .ZN(new_n654));
  INV_X1    g0454(.A(new_n643), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT92), .B1(new_n632), .B2(new_n639), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n632), .A2(new_n650), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n658), .A2(new_n651), .A3(new_n649), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n614), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n482), .A2(new_n545), .A3(new_n663), .ZN(G372));
  XNOR2_X1  g0464(.A(new_n384), .B(KEYINPUT98), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT18), .B1(new_n461), .B2(new_n472), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n458), .A2(new_n475), .A3(new_n474), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n460), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n392), .A2(new_n389), .A3(new_n388), .ZN(new_n671));
  INV_X1    g0471(.A(new_n373), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n341), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n669), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n296), .B1(new_n665), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n578), .B1(new_n560), .B2(new_n579), .ZN(new_n676));
  INV_X1    g0476(.A(new_n580), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n570), .A2(new_n573), .A3(new_n582), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n561), .B2(new_n574), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n644), .A2(new_n652), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n680), .A2(new_n681), .A3(new_n544), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n605), .A2(new_n610), .A3(new_n612), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n539), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n644), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n575), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n644), .A2(KEYINPUT93), .A3(new_n652), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n660), .B1(new_n657), .B2(new_n659), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT26), .B(new_n687), .C1(new_n688), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n687), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n675), .B1(new_n482), .B2(new_n696), .ZN(G369));
  NAND3_X1  g0497(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n704), .B1(new_n509), .B2(new_n516), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n545), .A2(new_n705), .B1(new_n539), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n603), .A2(new_n704), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n683), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n613), .B2(new_n707), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT99), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n534), .A2(new_n541), .A3(new_n544), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n684), .A2(new_n703), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n703), .B(KEYINPUT100), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n517), .A2(new_n533), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n712), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n207), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n627), .A2(G116), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n218), .B2(new_n722), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n713), .A2(new_n662), .A3(new_n614), .A4(new_n716), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n528), .A2(new_n621), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n609), .A3(new_n576), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(new_n609), .A3(new_n732), .A4(new_n576), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n606), .A2(new_n648), .A3(G179), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n532), .A3(new_n560), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n704), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n736), .ZN(new_n739));
  INV_X1    g0539(.A(new_n716), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT101), .B(KEYINPUT31), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n727), .B1(new_n728), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n662), .A2(new_n687), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT102), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(new_n692), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n575), .B1(new_n653), .B2(new_n661), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT102), .B1(new_n748), .B2(KEYINPUT26), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n747), .B(new_n749), .C1(new_n692), .C2(new_n691), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n534), .A2(new_n541), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n684), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n644), .B1(new_n752), .B2(new_n682), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n703), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT29), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n740), .B1(new_n686), .B2(new_n694), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT29), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n744), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n726), .B1(new_n758), .B2(G1), .ZN(G364));
  AND2_X1   g0559(.A1(new_n204), .A2(G13), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G45), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT103), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n763), .A2(new_n203), .A3(new_n721), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n710), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G330), .B2(new_n709), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n293), .A2(KEYINPUT105), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n204), .B1(KEYINPUT105), .B2(new_n293), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n210), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n579), .A2(new_n363), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n204), .A2(G179), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(G303), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n204), .A2(new_n370), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(new_n363), .A3(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G317), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(KEYINPUT33), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n776), .B(new_n784), .C1(G329), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n778), .A2(new_n579), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n772), .ZN(new_n792));
  INV_X1    g0592(.A(G326), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n773), .A2(new_n579), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n257), .B(new_n794), .C1(G283), .C2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n579), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n204), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G294), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT106), .ZN(new_n802));
  AND3_X1   g0602(.A1(new_n777), .A2(new_n802), .A3(new_n785), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n777), .B2(new_n785), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G311), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n788), .A2(new_n797), .A3(new_n801), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n795), .A2(new_n355), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n792), .A2(new_n222), .B1(new_n774), .B2(new_n491), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n809), .B(new_n810), .C1(new_n274), .C2(new_n789), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n799), .A2(new_n566), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n490), .B(new_n812), .C1(G68), .C2(new_n779), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n806), .A2(G77), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n786), .A2(new_n420), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT32), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n811), .A2(new_n813), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n771), .B1(new_n808), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G13), .A2(G33), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n204), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT104), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n771), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n219), .A2(new_n524), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n720), .A2(new_n408), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n823), .B(new_n824), .C1(new_n524), .C2(new_n248), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n720), .A2(new_n490), .ZN(new_n826));
  INV_X1    g0626(.A(G116), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n826), .A2(G355), .B1(new_n827), .B2(new_n720), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n764), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n818), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n709), .B2(new_n821), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n766), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n372), .A2(new_n703), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n368), .A2(new_n373), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT108), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n672), .A2(new_n703), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n368), .A2(new_n373), .A3(new_n835), .A4(KEYINPUT108), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n756), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT26), .B1(new_n681), .B2(new_n687), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n748), .B2(KEYINPUT26), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n680), .A2(new_n681), .A3(new_n544), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n683), .B1(new_n517), .B2(new_n533), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n657), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n716), .B(new_n841), .C1(new_n844), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT109), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n695), .A2(KEYINPUT109), .A3(new_n716), .A4(new_n841), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n852), .A2(new_n744), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n764), .B1(new_n852), .B2(new_n744), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(KEYINPUT110), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(KEYINPUT110), .B2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n792), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n779), .A2(G150), .B1(new_n857), .B2(G137), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n859), .B2(new_n790), .C1(new_n805), .C2(new_n420), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n774), .A2(new_n222), .B1(new_n786), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G68), .B2(new_n796), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n547), .B1(new_n800), .B2(new_n274), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n787), .A2(G311), .ZN(new_n867));
  INV_X1    g0667(.A(G283), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n780), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(G294), .B2(new_n789), .ZN(new_n870));
  INV_X1    g0670(.A(new_n812), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n792), .A2(new_n775), .B1(new_n774), .B2(new_n355), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n257), .B(new_n872), .C1(G87), .C2(new_n796), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n806), .A2(new_n500), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n771), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n770), .A2(new_n819), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT107), .Z(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n830), .B(new_n876), .C1(new_n224), .C2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n819), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n841), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n856), .A2(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n568), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n211), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(KEYINPUT111), .B(KEYINPUT36), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n216), .A2(G77), .A3(new_n217), .A4(new_n418), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n222), .A2(G68), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n203), .B(G13), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n701), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n669), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n428), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n441), .B1(new_n405), .B2(new_n411), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n457), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n701), .B1(new_n899), .B2(new_n446), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n473), .A2(new_n476), .A3(new_n477), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n479), .A2(new_n456), .A3(new_n459), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT112), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT112), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n480), .A2(new_n905), .A3(new_n900), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n461), .B1(new_n472), .B2(new_n894), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n454), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n899), .A2(new_n446), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n472), .B2(new_n894), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .A3(new_n454), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n903), .A2(KEYINPUT112), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n905), .B1(new_n480), .B2(new_n900), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT113), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n917), .B1(new_n904), .B2(new_n906), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT113), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n916), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n373), .A2(new_n703), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT109), .B1(new_n756), .B2(new_n841), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n848), .A2(new_n849), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n317), .A2(new_n703), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n340), .A2(new_n671), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n334), .A2(G169), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT14), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n337), .A3(new_n336), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n391), .B2(new_n393), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n931), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n896), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n341), .A2(new_n704), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n456), .B(new_n459), .C1(new_n666), .C2(new_n667), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n458), .A2(new_n701), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n458), .B1(new_n475), .B2(new_n701), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT37), .B1(new_n945), .B2(KEYINPUT114), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n943), .A2(new_n944), .B1(new_n946), .B2(new_n909), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n909), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT39), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n926), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n940), .B1(new_n942), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n755), .A2(new_n481), .A3(new_n757), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n955), .A2(new_n675), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n737), .B2(new_n741), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n728), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n936), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n932), .B1(new_n394), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n340), .A2(new_n671), .A3(new_n932), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n841), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n958), .B1(new_n926), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n958), .B(new_n967), .C1(new_n728), .C2(new_n961), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n924), .B2(new_n949), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT115), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n971), .B(KEYINPUT115), .C1(new_n924), .C2(new_n949), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n970), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n482), .B2(new_n963), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n970), .A2(new_n481), .A3(new_n962), .A4(new_n976), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(G330), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n957), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n203), .B2(new_n760), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n957), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n893), .B1(new_n982), .B2(new_n983), .ZN(G367));
  INV_X1    g0784(.A(new_n822), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n207), .B2(new_n346), .ZN(new_n986));
  INV_X1    g0786(.A(new_n824), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n244), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n764), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n795), .A2(new_n566), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n787), .ZN(new_n991));
  INV_X1    g0791(.A(new_n774), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  INV_X1    g0793(.A(G294), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n993), .C1(new_n994), .C2(new_n780), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G283), .B2(new_n806), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n789), .A2(G303), .B1(new_n857), .B2(G311), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT119), .Z(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT46), .B1(new_n992), .B2(new_n500), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n408), .B(new_n999), .C1(new_n359), .C2(new_n800), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n796), .A2(G77), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n859), .B2(new_n792), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n490), .B(new_n1003), .C1(G137), .C2(new_n787), .ZN(new_n1004));
  INV_X1    g0804(.A(G150), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1005), .A2(new_n790), .B1(new_n780), .B2(new_n420), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n274), .B2(new_n992), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n800), .A2(G68), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n806), .A2(G50), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n989), .B1(new_n1012), .B2(new_n770), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n658), .A2(new_n704), .ZN(new_n1014));
  MUX2_X1   g0814(.A(new_n681), .B(new_n644), .S(new_n1014), .Z(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1015), .B2(new_n821), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n763), .A2(new_n203), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n574), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n680), .B1(new_n1019), .B2(new_n716), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n687), .A2(new_n740), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n718), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT45), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(KEYINPUT118), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n718), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1026), .A2(KEYINPUT118), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n712), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n715), .B1(new_n706), .B2(new_n714), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(new_n710), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n758), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n758), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n721), .B(KEYINPUT41), .Z(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1018), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT117), .Z(new_n1041));
  NAND3_X1  g0841(.A1(new_n713), .A2(new_n1022), .A3(new_n714), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT42), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT42), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n575), .B1(new_n751), .B2(new_n1020), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n716), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1041), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT116), .Z(new_n1050));
  XNOR2_X1  g0850(.A(new_n1048), .B(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n712), .A2(new_n1022), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1051), .B(new_n1052), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n1016), .B1(new_n1039), .B2(new_n1053), .ZN(G387));
  OR2_X1    g0854(.A1(new_n706), .A2(new_n821), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n824), .B1(new_n241), .B2(new_n524), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n826), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n723), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n343), .A2(new_n222), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT50), .Z(new_n1060));
  AOI21_X1  g0860(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n723), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1058), .A2(new_n1062), .B1(new_n355), .B2(new_n720), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n764), .B1(new_n1063), .B2(new_n822), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n789), .A2(G50), .B1(new_n857), .B2(G159), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1005), .B2(new_n786), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n774), .A2(new_n224), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1066), .A2(new_n547), .A3(new_n990), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n806), .A2(G68), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n779), .A2(new_n275), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n637), .A2(new_n800), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G311), .A2(new_n779), .B1(new_n789), .B2(G317), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n791), .B2(new_n792), .C1(new_n805), .C2(new_n775), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n800), .A2(G283), .B1(new_n992), .B2(G294), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n795), .A2(new_n499), .B1(new_n786), .B2(new_n793), .ZN(new_n1082));
  OR3_X1    g0882(.A1(new_n1081), .A2(new_n408), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1072), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1064), .B1(new_n1085), .B2(new_n770), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1034), .A2(new_n1018), .B1(new_n1055), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1035), .A2(new_n721), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n758), .A2(new_n1034), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT120), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(G393));
  AND2_X1   g0894(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n721), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1032), .A2(new_n1017), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n985), .B1(new_n566), .B2(new_n207), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n987), .A2(new_n251), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n764), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n789), .A2(G311), .B1(new_n857), .B2(G317), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n806), .A2(G294), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n780), .A2(new_n775), .B1(new_n786), .B2(new_n791), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G283), .B2(new_n992), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n257), .B(new_n809), .C1(new_n500), .C2(new_n800), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n789), .A2(G159), .B1(new_n857), .B2(G150), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT51), .Z(new_n1110));
  OAI22_X1  g0910(.A1(new_n795), .A2(new_n491), .B1(new_n786), .B2(new_n859), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n227), .B2(new_n992), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n800), .A2(G77), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1110), .A2(new_n408), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n806), .A2(new_n343), .B1(G50), .B2(new_n779), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT121), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1108), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1101), .B1(new_n1117), .B2(new_n770), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1022), .B2(new_n821), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1098), .A2(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1097), .A2(new_n1120), .ZN(G390));
  AOI21_X1  g0921(.A(new_n927), .B1(new_n850), .B2(new_n851), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n938), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n941), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n951), .B(new_n1124), .C1(new_n926), .C2(new_n952), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n947), .A2(new_n948), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT38), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n921), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n838), .A2(new_n840), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n927), .B1(new_n754), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n938), .B(KEYINPUT122), .Z(new_n1132));
  OAI211_X1 g0932(.A(new_n941), .B(new_n1129), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n841), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n727), .B(new_n1134), .C1(new_n728), .C2(new_n743), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n938), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1125), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n750), .A2(new_n753), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n704), .A3(new_n1130), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1132), .B1(new_n1139), .B2(new_n928), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1129), .A2(new_n941), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1127), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT113), .B1(new_n907), .B2(new_n918), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n922), .B(new_n917), .C1(new_n904), .C2(new_n906), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n950), .B1(new_n1147), .B2(KEYINPUT39), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1148), .B2(new_n1124), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1134), .A2(new_n727), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n962), .A2(new_n938), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1137), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n481), .A2(new_n962), .A3(G330), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT123), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n955), .A3(new_n675), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n962), .A2(new_n1150), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1135), .A2(new_n938), .B1(new_n1156), .B2(new_n1132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1135), .B2(new_n938), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1131), .A2(new_n1157), .B1(new_n931), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1152), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1137), .B(new_n1160), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n721), .A3(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1137), .B(new_n1018), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n764), .B1(new_n878), .B2(new_n275), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n774), .A2(new_n1005), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT53), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n257), .B1(new_n1167), .B2(new_n792), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n789), .A2(G132), .B1(G50), .B2(new_n796), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n786), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1170), .B(new_n1173), .C1(new_n1169), .C2(new_n1168), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G137), .A2(new_n779), .B1(new_n800), .B2(G159), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n805), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT124), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n779), .A2(new_n359), .B1(new_n857), .B2(G283), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n994), .B2(new_n786), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G97), .B2(new_n806), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n257), .B1(new_n992), .B2(G87), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n789), .A2(G116), .B1(G68), .B2(new_n796), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n1113), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1179), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1186), .B2(new_n770), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n953), .B2(new_n881), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1165), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1164), .A2(new_n1189), .ZN(G378));
  INV_X1    g0990(.A(KEYINPUT125), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n895), .B1(new_n1147), .B2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n1148), .B2(new_n941), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n727), .B1(new_n974), .B2(new_n975), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n665), .A2(new_n295), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n292), .A2(new_n894), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1199), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1196), .B1(new_n292), .B2(new_n894), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n665), .B2(new_n295), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n970), .A2(new_n1195), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n970), .B2(new_n1195), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1194), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n970), .A2(new_n1195), .A3(new_n1205), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT115), .B1(new_n1129), .B2(new_n971), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n967), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n663), .A2(new_n545), .A3(new_n740), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(KEYINPUT40), .C1(new_n1213), .C2(new_n960), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n973), .B(new_n1214), .C1(new_n921), .C2(new_n1128), .ZN(new_n1215));
  OAI21_X1  g1015(.A(G330), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT40), .B1(new_n1147), .B2(new_n968), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n954), .A2(new_n1209), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1017), .B1(new_n1208), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1205), .A2(new_n881), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n408), .A2(G41), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n796), .A2(new_n274), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1008), .B(new_n1225), .C1(new_n224), .C2(new_n774), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n780), .A2(new_n566), .B1(new_n792), .B2(new_n827), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n790), .A2(new_n355), .B1(new_n786), .B2(new_n868), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n1222), .C1(new_n634), .C2(new_n805), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1224), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n792), .A2(new_n1172), .B1(new_n774), .B2(new_n1176), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1167), .A2(new_n790), .B1(new_n780), .B2(new_n862), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(G150), .C2(new_n800), .ZN(new_n1235));
  INV_X1    g1035(.A(G137), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n805), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n796), .A2(G159), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n770), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n764), .C1(G50), .C2(new_n878), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1221), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1191), .B1(new_n1220), .B2(new_n1246), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1206), .A2(new_n1207), .A3(new_n1194), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n953), .A2(new_n942), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1218), .A2(new_n1209), .B1(new_n1249), .B2(new_n1193), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1018), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1246), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(KEYINPUT125), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1247), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1208), .A2(new_n1219), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1155), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1163), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1257), .A3(KEYINPUT57), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1219), .A2(new_n1208), .B1(new_n1163), .B2(new_n1256), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n721), .C1(KEYINPUT57), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(G375));
  INV_X1    g1061(.A(new_n1159), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1132), .A2(new_n819), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n764), .B1(new_n878), .B2(G68), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n790), .A2(new_n868), .B1(new_n792), .B2(new_n994), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G303), .B2(new_n787), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n779), .A2(new_n500), .B1(G97), .B2(new_n992), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1266), .A2(new_n490), .A3(new_n1002), .A4(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1071), .B1(new_n496), .B2(new_n805), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n800), .A2(G50), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n787), .A2(G128), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n408), .A3(new_n1225), .A4(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1176), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n779), .A2(new_n1273), .B1(new_n857), .B2(G132), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n789), .A2(G137), .B1(G159), .B2(new_n992), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(new_n805), .C2(new_n1005), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1268), .A2(new_n1269), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1264), .B1(new_n1277), .B2(new_n770), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1262), .A2(new_n1018), .B1(new_n1263), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1161), .A2(new_n1038), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(G381));
  AND2_X1   g1082(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1283));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(G390), .A2(G387), .A3(G384), .A4(G381), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(G407));
  NAND2_X1  g1087(.A1(new_n702), .A2(G213), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G407), .B(G213), .C1(G375), .C2(new_n1290), .ZN(G409));
  INV_X1    g1091(.A(KEYINPUT127), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(G393), .B(new_n833), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1097), .A2(new_n1120), .ZN(new_n1294));
  AND2_X1   g1094(.A1(G387), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1293), .B1(new_n1295), .B2(KEYINPUT126), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G387), .A2(new_n1294), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(new_n1294), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1293), .A3(KEYINPUT126), .A4(new_n1298), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1254), .A2(new_n1260), .A3(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1259), .A2(new_n1038), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1284), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1289), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1281), .A2(new_n1309), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1256), .A2(new_n1262), .A3(KEYINPUT60), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n721), .B(new_n1161), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1312), .B2(new_n1279), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(G384), .A3(new_n1279), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1289), .A2(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1314), .A2(new_n1315), .A3(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1303), .B1(new_n1308), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1316), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1308), .B2(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1322), .A2(new_n1325), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1289), .B(new_n1316), .C1(new_n1304), .C2(new_n1307), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1323), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1302), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1308), .A2(KEYINPUT63), .A3(new_n1324), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1330), .B(new_n1303), .C1(new_n1308), .C2(new_n1321), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1302), .B1(new_n1327), .B2(KEYINPUT63), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1292), .B1(new_n1329), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1322), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1308), .A2(new_n1324), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1335), .A2(new_n1338), .A3(new_n1302), .A4(new_n1330), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1340), .A2(new_n1322), .A3(new_n1325), .ZN(new_n1341));
  OAI211_X1 g1141(.A(KEYINPUT127), .B(new_n1339), .C1(new_n1341), .C2(new_n1302), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1334), .A2(new_n1342), .ZN(G405));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1284), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1304), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1316), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1302), .ZN(G402));
endmodule


