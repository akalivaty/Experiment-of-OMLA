//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204));
  AND3_X1   g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT2), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n203), .B2(KEYINPUT2), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  INV_X1    g008(.A(G141gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT79), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n203), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n207), .A2(new_n212), .A3(new_n215), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT78), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n225), .A3(KEYINPUT2), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n212), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n213), .A2(new_n214), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND4_X1   g028(.A1(new_n202), .A2(new_n221), .A3(new_n222), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n229), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT81), .B1(new_n232), .B2(KEYINPUT3), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G211gat), .B(G218gat), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G211gat), .A2(G218gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(KEYINPUT72), .B2(KEYINPUT22), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT73), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT72), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT22), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n242), .A2(new_n243), .B1(G211gat), .B2(G218gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n239), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G197gat), .B(G204gat), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n236), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  AOI211_X1 g049(.A(new_n235), .B(new_n248), .C1(new_n241), .C2(new_n246), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n215), .A2(new_n220), .A3(new_n212), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n255), .A2(new_n207), .B1(new_n228), .B2(new_n227), .ZN(new_n256));
  INV_X1    g055(.A(new_n250), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n247), .A2(new_n236), .A3(new_n249), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT88), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT29), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n250), .B2(new_n251), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT3), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n256), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G228gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  OAI22_X1  g066(.A1(new_n254), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n266), .B(new_n267), .C1(new_n259), .C2(new_n232), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n232), .A2(KEYINPUT3), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n269), .B(new_n270), .C1(new_n253), .C2(new_n234), .ZN(new_n271));
  XOR2_X1   g070(.A(G78gat), .B(G106gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT31), .ZN(new_n273));
  INV_X1    g072(.A(G50gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n268), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G22gat), .ZN(new_n278));
  INV_X1    g077(.A(G22gat), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n268), .A2(new_n279), .A3(new_n271), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n268), .A2(new_n271), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT89), .B1(new_n282), .B2(new_n275), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n281), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G120gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT1), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G127gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n295), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n287), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  OAI21_X1  g097(.A(G127gat), .B1(new_n295), .B2(KEYINPUT1), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(G134gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n302), .B1(KEYINPUT26), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n304), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT28), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n320), .A3(new_n317), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  AND2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n305), .A3(new_n306), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n323), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n302), .B2(KEYINPUT24), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n302), .B2(KEYINPUT24), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT66), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n328), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n328), .B2(new_n335), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n327), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n309), .ZN(new_n342));
  AOI211_X1 g141(.A(KEYINPUT65), .B(new_n324), .C1(new_n326), .C2(new_n327), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n333), .A2(KEYINPUT64), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n330), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n301), .B(new_n322), .C1(new_n339), .C2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n297), .A2(new_n300), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n335), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT67), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n328), .A2(new_n335), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n341), .A2(new_n309), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT65), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n340), .A3(new_n309), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n347), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n354), .A2(new_n355), .B1(new_n359), .B2(new_n323), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n319), .A2(new_n321), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n314), .B2(new_n312), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n354), .A2(new_n355), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n323), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(KEYINPUT69), .A3(new_n301), .A4(new_n322), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n286), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT33), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n370), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  AOI221_X4 g175(.A(new_n286), .B1(KEYINPUT33), .B2(new_n374), .C1(new_n368), .C2(new_n369), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n285), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n368), .A2(new_n369), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT70), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n368), .A2(new_n369), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT33), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n370), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n377), .ZN(new_n387));
  INV_X1    g186(.A(new_n285), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n378), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n381), .B1(new_n378), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n284), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n297), .A2(new_n229), .A3(new_n221), .A4(new_n300), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n256), .A2(new_n395), .A3(new_n300), .A4(new_n297), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(KEYINPUT86), .A3(new_n396), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n393), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n232), .A2(KEYINPUT3), .B1(new_n297), .B2(new_n300), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n202), .B1(new_n256), .B2(new_n222), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n230), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT5), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(KEYINPUT82), .A3(new_n396), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n408), .A3(KEYINPUT4), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n407), .A2(new_n402), .A3(new_n404), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n352), .A2(new_n232), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n393), .ZN(new_n412));
  INV_X1    g211(.A(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n410), .A2(KEYINPUT83), .A3(new_n414), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n406), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT85), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT87), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT6), .B1(new_n419), .B2(new_n425), .ZN(new_n427));
  INV_X1    g226(.A(new_n418), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT83), .B1(new_n410), .B2(new_n414), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n428), .A2(new_n429), .B1(new_n399), .B2(new_n405), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G8gat), .B(G36gat), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G64gat), .ZN(new_n438));
  INV_X1    g237(.A(G92gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n442));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n442), .B2(KEYINPUT29), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(KEYINPUT74), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n442), .A2(new_n447), .A3(new_n443), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n446), .A2(new_n253), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT75), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n444), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n261), .B1(new_n360), .B2(new_n362), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT75), .A3(new_n443), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n252), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT30), .B(new_n441), .C1(new_n449), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n451), .A2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n253), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n440), .B(KEYINPUT76), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n448), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n447), .B1(new_n452), .B2(new_n443), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n252), .C1(new_n462), .C2(new_n444), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n455), .A2(new_n456), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n463), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT30), .B1(new_n467), .B2(new_n441), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n455), .A2(new_n464), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT77), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n436), .A2(new_n466), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n392), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n449), .A2(new_n454), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n440), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n464), .A3(new_n455), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n427), .B1(new_n425), .B2(new_n419), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n476), .B1(new_n435), .B2(new_n477), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n376), .A2(new_n285), .A3(new_n377), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n388), .B1(new_n386), .B2(new_n387), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n380), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n378), .A2(new_n381), .A3(new_n389), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n478), .A2(new_n483), .A3(new_n484), .A4(new_n284), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n472), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n284), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n413), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n425), .B1(new_n490), .B2(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n411), .A2(new_n404), .A3(new_n393), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT39), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT90), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n495), .A2(KEYINPUT40), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n495), .A2(KEYINPUT40), .B1(new_n430), .B2(new_n432), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(new_n497), .C1(new_n469), .C2(new_n468), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n458), .A2(new_n499), .A3(new_n463), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n457), .A2(new_n252), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n461), .B(new_n253), .C1(new_n462), .C2(new_n444), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT37), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n459), .A2(KEYINPUT38), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n477), .A2(new_n506), .A3(new_n435), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT37), .B1(new_n449), .B2(new_n454), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n441), .B1(new_n500), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT38), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n509), .A2(new_n510), .B1(new_n474), .B2(new_n440), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n284), .B(new_n498), .C1(new_n507), .C2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n481), .A2(KEYINPUT36), .A3(new_n482), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n390), .B2(new_n391), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n488), .A2(new_n512), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518));
  XNOR2_X1  g317(.A(G183gat), .B(G211gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G15gat), .B(G22gat), .Z(new_n522));
  OR2_X1    g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  INV_X1    g322(.A(G1gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G8gat), .ZN(new_n530));
  INV_X1    g329(.A(G8gat), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n523), .A2(new_n526), .A3(new_n531), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT21), .ZN(new_n535));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538));
  INV_X1    g337(.A(G71gat), .ZN(new_n539));
  INV_X1    g338(.A(G78gat), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G57gat), .B(G64gat), .Z(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n534), .B1(new_n535), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT95), .ZN(new_n548));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n549), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n521), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(new_n521), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n546), .A2(new_n535), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n553), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n553), .B2(new_n556), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n439), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n565), .B2(new_n439), .ZN(new_n568));
  NAND3_X1  g367(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n570), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n576));
  INV_X1    g375(.A(G29gat), .ZN(new_n577));
  INV_X1    g376(.A(G36gat), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n579), .B2(KEYINPUT91), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n581));
  NOR2_X1   g380(.A1(G29gat), .A2(G36gat), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n576), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n574), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G43gat), .B(G50gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT15), .A3(new_n585), .ZN(new_n586));
  OR3_X1    g385(.A1(new_n585), .A2(KEYINPUT92), .A3(KEYINPUT15), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n585), .B2(KEYINPUT15), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n585), .A2(KEYINPUT15), .B1(new_n579), .B2(new_n575), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n587), .A2(new_n574), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT17), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n586), .B2(new_n590), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n573), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n570), .B(new_n571), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G190gat), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n595), .A2(new_n317), .A3(new_n596), .A4(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G218gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(G218gat), .A3(new_n601), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT96), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT97), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n608), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n604), .A2(new_n614), .A3(new_n605), .A4(new_n609), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n563), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n545), .A3(new_n543), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n573), .A2(new_n546), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n545), .A4(new_n543), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n619), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n306), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G204gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n629), .A2(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n518), .B1(new_n617), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n562), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n637), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(KEYINPUT98), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n517), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n534), .B1(new_n592), .B2(new_n594), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT94), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n533), .A2(new_n591), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n534), .B(new_n648), .C1(new_n592), .C2(new_n594), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n533), .B(new_n591), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n647), .B(KEYINPUT13), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT11), .B(G169gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G197gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G113gat), .B(G141gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT12), .Z(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n650), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n650), .A2(new_n663), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n664), .A2(new_n660), .A3(new_n654), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n643), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n436), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n524), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT42), .ZN(new_n671));
  INV_X1    g470(.A(new_n668), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n476), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n673), .B2(G8gat), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n476), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(KEYINPUT99), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(KEYINPUT99), .B2(KEYINPUT42), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n674), .A2(new_n676), .B1(new_n678), .B2(new_n679), .ZN(G1325gat));
  AOI21_X1  g479(.A(G15gat), .B1(new_n672), .B2(new_n483), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n668), .B1(new_n513), .B2(new_n515), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n681), .B1(G15gat), .B2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n284), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n517), .B2(new_n639), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n688), .B(new_n616), .C1(new_n486), .C2(new_n516), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n691));
  INV_X1    g490(.A(new_n436), .ZN(new_n692));
  INV_X1    g491(.A(new_n667), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n563), .A2(new_n693), .A3(new_n637), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n690), .A2(new_n691), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n515), .A2(new_n513), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n465), .B1(new_n434), .B2(new_n435), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n284), .B1(new_n697), .B2(new_n470), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n699), .A2(new_n512), .B1(new_n472), .B2(new_n485), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n688), .B1(new_n700), .B2(new_n616), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n517), .A2(KEYINPUT44), .A3(new_n639), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n701), .A2(new_n692), .A3(new_n702), .A4(new_n694), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n695), .A2(new_n704), .A3(G29gat), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n517), .A2(new_n639), .A3(new_n694), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n577), .A3(new_n692), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n706), .A2(new_n709), .A3(new_n577), .A4(new_n692), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT101), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n705), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n706), .A2(new_n578), .A3(new_n476), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT46), .Z(new_n718));
  AND3_X1   g517(.A1(new_n690), .A2(new_n476), .A3(new_n694), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n578), .B2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n701), .A2(new_n696), .A3(new_n702), .A4(new_n694), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n721), .A3(new_n483), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(KEYINPUT47), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(G43gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n726), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n727), .A2(new_n731), .ZN(G1330gat));
  NAND3_X1  g531(.A1(new_n690), .A2(new_n487), .A3(new_n694), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT48), .B1(new_n734), .B2(KEYINPUT104), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n706), .A2(new_n274), .A3(new_n487), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(new_n736), .C1(KEYINPUT104), .C2(KEYINPUT48), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1331gat));
  NOR4_X1   g539(.A1(new_n700), .A2(new_n667), .A3(new_n617), .A4(new_n641), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n692), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n476), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT49), .B(G64gat), .Z(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(G1333gat));
  XNOR2_X1  g546(.A(new_n483), .B(KEYINPUT105), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n741), .A2(new_n539), .A3(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n741), .A2(new_n696), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n539), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g551(.A1(new_n741), .A2(new_n487), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n563), .A2(new_n667), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n517), .A2(new_n639), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT106), .B(KEYINPUT51), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(KEYINPUT106), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n692), .A2(new_n565), .A3(new_n637), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT107), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n755), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n641), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n690), .A2(new_n692), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n565), .ZN(G1336gat));
  NAND3_X1  g568(.A1(new_n690), .A2(new_n476), .A3(new_n767), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n760), .B1(new_n757), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n756), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n476), .A2(new_n439), .A3(new_n637), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n780), .A3(new_n776), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n771), .A3(new_n779), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n762), .B2(new_n776), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n778), .A2(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1337gat));
  AOI21_X1  g583(.A(new_n641), .B1(new_n759), .B2(new_n761), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT110), .B(G99gat), .Z(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n483), .A3(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n690), .A2(new_n696), .A3(new_n767), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(G1338gat));
  NOR2_X1   g589(.A1(new_n284), .A2(G106gat), .ZN(new_n791));
  AND4_X1   g590(.A1(new_n637), .A2(new_n773), .A3(new_n774), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n690), .A2(new_n487), .A3(new_n767), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT53), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT53), .B1(new_n785), .B2(new_n791), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n793), .A2(KEYINPUT111), .ZN(new_n797));
  OAI21_X1  g596(.A(G106gat), .B1(new_n793), .B2(KEYINPUT111), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(G1339gat));
  NAND3_X1  g599(.A1(new_n621), .A2(new_n622), .A3(new_n627), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n625), .A2(new_n801), .A3(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n627), .B1(new_n621), .B2(new_n622), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n632), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n802), .A2(KEYINPUT55), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT55), .B1(new_n802), .B2(new_n805), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n634), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n662), .B2(new_n666), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n811));
  INV_X1    g610(.A(new_n647), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n811), .A2(KEYINPUT112), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT112), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n652), .A2(new_n653), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n666), .B(new_n637), .C1(new_n816), .C2(new_n659), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n616), .B1(new_n810), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n808), .B(new_n666), .C1(new_n816), .C2(new_n659), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT113), .B1(new_n616), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n820), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n639), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n819), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n819), .A2(new_n821), .A3(new_n827), .A4(new_n824), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n562), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n640), .A2(new_n693), .A3(new_n641), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n392), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n476), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n692), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n667), .A2(new_n290), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT116), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n839), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n693), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n290), .ZN(G1340gat));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n288), .A3(new_n637), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n641), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n288), .ZN(G1341gat));
  AOI21_X1  g645(.A(G127gat), .B1(new_n835), .B2(new_n563), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n562), .B1(new_n840), .B2(new_n841), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(G127gat), .ZN(G1342gat));
  NAND3_X1  g648(.A1(new_n835), .A2(new_n287), .A3(new_n639), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n616), .B1(new_n840), .B2(new_n841), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n287), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n696), .A2(new_n833), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n821), .A2(new_n824), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n660), .B1(new_n651), .B2(new_n654), .ZN(new_n859));
  INV_X1    g658(.A(new_n666), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n639), .B1(new_n861), .B2(new_n817), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n562), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n830), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n487), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT118), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n867), .A3(KEYINPUT57), .A4(new_n487), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n284), .B1(new_n829), .B2(new_n830), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n667), .B(new_n855), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n829), .A2(new_n830), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n210), .A3(new_n487), .A4(new_n855), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n693), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT58), .B1(new_n876), .B2(KEYINPUT120), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(KEYINPUT120), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT119), .B1(new_n875), .B2(new_n693), .ZN(new_n880));
  INV_X1    g679(.A(new_n855), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n284), .B(new_n881), .C1(new_n829), .C2(new_n830), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n210), .A4(new_n667), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(G141gat), .B2(new_n872), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(G1344gat));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n870), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n638), .A2(new_n693), .A3(new_n642), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n862), .B1(new_n639), .B2(new_n822), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n563), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n889), .B(new_n487), .C1(new_n891), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n890), .A2(new_n637), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n855), .B(KEYINPUT121), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT59), .B(G148gat), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n208), .A3(new_n637), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n637), .B(new_n855), .C1(new_n869), .C2(new_n871), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(G148gat), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n897), .B(new_n898), .C1(new_n900), .C2(KEYINPUT59), .ZN(G1345gat));
  OR2_X1    g700(.A1(new_n869), .A2(new_n871), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n902), .A2(G155gat), .A3(new_n563), .A4(new_n855), .ZN(new_n903));
  INV_X1    g702(.A(new_n882), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n216), .B1(new_n904), .B2(new_n562), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(G1346gat));
  NAND4_X1  g705(.A1(new_n902), .A2(G162gat), .A3(new_n639), .A4(new_n855), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n217), .B1(new_n904), .B2(new_n616), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n692), .A2(new_n832), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n831), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n305), .A3(new_n667), .ZN(new_n912));
  INV_X1    g711(.A(new_n910), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n487), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n874), .A2(new_n748), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n693), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(G1348gat));
  NOR3_X1   g718(.A1(new_n915), .A2(new_n306), .A3(new_n641), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n911), .A2(new_n637), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n306), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n911), .A2(new_n563), .A3(new_n316), .ZN(new_n923));
  OAI21_X1  g722(.A(G183gat), .B1(new_n915), .B2(new_n562), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g725(.A1(new_n874), .A2(new_n639), .A3(new_n748), .A4(new_n914), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G190gat), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(KEYINPUT61), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n317), .A3(new_n639), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n913), .A2(new_n696), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n890), .A2(new_n894), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n693), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n870), .A2(new_n937), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(G197gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n693), .B2(new_n941), .ZN(G1352gat));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n870), .A2(new_n943), .A3(new_n637), .A4(new_n937), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  INV_X1    g745(.A(new_n937), .ZN(new_n947));
  OAI21_X1  g746(.A(G204gat), .B1(new_n895), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT124), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(G1353gat));
  OR3_X1    g750(.A1(new_n940), .A2(G211gat), .A3(new_n562), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n890), .A2(new_n563), .A3(new_n894), .A4(new_n937), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(new_n603), .B1(new_n940), .B2(new_n616), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n960));
  INV_X1    g759(.A(new_n938), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n639), .A2(G218gat), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT127), .Z(new_n963));
  AOI22_X1  g762(.A1(new_n959), .A2(new_n960), .B1(new_n961), .B2(new_n963), .ZN(G1355gat));
endmodule


