

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761;

  AND2_X1 U381 ( .A1(n680), .A2(n681), .ZN(n418) );
  AND2_X1 U382 ( .A1(n641), .A2(KEYINPUT44), .ZN(n379) );
  OR2_X1 U383 ( .A1(n646), .A2(n645), .ZN(n442) );
  NOR2_X2 U384 ( .A1(G953), .A2(G237), .ZN(n526) );
  XNOR2_X1 U385 ( .A(n393), .B(n477), .ZN(n478) );
  OR2_X1 U386 ( .A1(n633), .A2(n659), .ZN(n588) );
  INV_X1 U387 ( .A(G953), .ZN(n753) );
  NOR2_X1 U388 ( .A1(n689), .A2(n678), .ZN(n482) );
  BUF_X2 U389 ( .A(n603), .Z(n359) );
  NOR2_X1 U390 ( .A1(n761), .A2(n759), .ZN(n422) );
  OR2_X1 U391 ( .A1(n435), .A2(n432), .ZN(n431) );
  NAND2_X1 U392 ( .A1(n608), .A2(n607), .ZN(n609) );
  INV_X1 U393 ( .A(KEYINPUT22), .ZN(n403) );
  NAND2_X1 U394 ( .A1(n634), .A2(n420), .ZN(n419) );
  XNOR2_X1 U395 ( .A(n611), .B(n459), .ZN(n626) );
  NAND2_X1 U396 ( .A1(n596), .A2(n590), .ZN(n611) );
  XNOR2_X1 U397 ( .A(n535), .B(n446), .ZN(n740) );
  XNOR2_X1 U398 ( .A(n741), .B(n412), .ZN(n393) );
  XNOR2_X1 U399 ( .A(n474), .B(n473), .ZN(n741) );
  XNOR2_X1 U400 ( .A(n465), .B(n464), .ZN(n535) );
  XNOR2_X1 U401 ( .A(G146), .B(G125), .ZN(n380) );
  NOR2_X2 U402 ( .A1(n396), .A2(n395), .ZN(n703) );
  NOR2_X2 U403 ( .A1(n758), .A2(n703), .ZN(n414) );
  NOR2_X1 U404 ( .A1(n694), .A2(G902), .ZN(n538) );
  XNOR2_X1 U405 ( .A(n525), .B(n524), .ZN(n541) );
  XNOR2_X1 U406 ( .A(G131), .B(G134), .ZN(n524) );
  XNOR2_X1 U407 ( .A(n541), .B(n361), .ZN(n748) );
  NAND2_X1 U408 ( .A1(n431), .A2(n439), .ZN(n673) );
  XNOR2_X1 U409 ( .A(G104), .B(G122), .ZN(n503) );
  INV_X1 U410 ( .A(KEYINPUT100), .ZN(n387) );
  XNOR2_X1 U411 ( .A(n380), .B(KEYINPUT10), .ZN(n747) );
  XNOR2_X1 U412 ( .A(G113), .B(G143), .ZN(n497) );
  XOR2_X1 U413 ( .A(G140), .B(G131), .Z(n498) );
  XOR2_X1 U414 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n501) );
  NAND2_X1 U415 ( .A1(n495), .A2(n458), .ZN(n457) );
  XNOR2_X1 U416 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n458) );
  NOR2_X1 U417 ( .A1(n618), .A2(n433), .ZN(n432) );
  NAND2_X1 U418 ( .A1(n619), .A2(n438), .ZN(n436) );
  XNOR2_X1 U419 ( .A(n382), .B(n381), .ZN(n610) );
  INV_X1 U420 ( .A(KEYINPUT108), .ZN(n381) );
  NAND2_X1 U421 ( .A1(n383), .A2(n712), .ZN(n382) );
  NOR2_X1 U422 ( .A1(n635), .A2(n384), .ZN(n383) );
  OR2_X1 U423 ( .A1(G237), .A2(G902), .ZN(n483) );
  XOR2_X1 U424 ( .A(KEYINPUT73), .B(G137), .Z(n531) );
  XNOR2_X1 U425 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n530) );
  XOR2_X1 U426 ( .A(G146), .B(KEYINPUT97), .Z(n528) );
  NOR2_X1 U427 ( .A1(n637), .A2(KEYINPUT106), .ZN(n399) );
  XNOR2_X1 U428 ( .A(n372), .B(n519), .ZN(n659) );
  OR2_X1 U429 ( .A1(n731), .A2(G902), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n731) );
  XNOR2_X1 U431 ( .A(n360), .B(n513), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n514), .B(n518), .ZN(n374) );
  XNOR2_X1 U433 ( .A(G119), .B(G110), .ZN(n513) );
  AND2_X1 U434 ( .A1(n681), .A2(G475), .ZN(n413) );
  XNOR2_X1 U435 ( .A(n440), .B(n748), .ZN(n725) );
  XNOR2_X1 U436 ( .A(n460), .B(n542), .ZN(n441) );
  INV_X1 U437 ( .A(G146), .ZN(n542) );
  XNOR2_X1 U438 ( .A(n690), .B(KEYINPUT54), .ZN(n691) );
  NAND2_X1 U439 ( .A1(n389), .A2(n388), .ZN(n439) );
  XNOR2_X1 U440 ( .A(n391), .B(n390), .ZN(n389) );
  INV_X1 U441 ( .A(KEYINPUT43), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n423), .B(n606), .ZN(n761) );
  INV_X1 U443 ( .A(KEYINPUT44), .ZN(n369) );
  INV_X1 U444 ( .A(KEYINPUT4), .ZN(n476) );
  INV_X1 U445 ( .A(KEYINPUT65), .ZN(n456) );
  NAND2_X1 U446 ( .A1(n434), .A2(KEYINPUT48), .ZN(n433) );
  INV_X1 U447 ( .A(n619), .ZN(n434) );
  XNOR2_X1 U448 ( .A(G902), .B(KEYINPUT15), .ZN(n480) );
  XNOR2_X1 U449 ( .A(G116), .B(G113), .ZN(n463) );
  XNOR2_X1 U450 ( .A(G110), .B(G104), .ZN(n472) );
  XNOR2_X1 U451 ( .A(n378), .B(KEYINPUT105), .ZN(n376) );
  NAND2_X1 U452 ( .A1(n444), .A2(n696), .ZN(n378) );
  XNOR2_X1 U453 ( .A(n421), .B(n467), .ZN(n469) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n467) );
  NAND2_X1 U455 ( .A1(G234), .A2(G237), .ZN(n566) );
  NOR2_X1 U456 ( .A1(n559), .A2(n635), .ZN(n560) );
  INV_X1 U457 ( .A(G469), .ZN(n454) );
  OR2_X1 U458 ( .A1(n725), .A2(G902), .ZN(n455) );
  XNOR2_X1 U459 ( .A(n649), .B(n443), .ZN(n646) );
  INV_X1 U460 ( .A(KEYINPUT93), .ZN(n443) );
  INV_X1 U461 ( .A(n633), .ZN(n420) );
  NAND2_X1 U462 ( .A1(n431), .A2(n363), .ZN(n751) );
  XOR2_X1 U463 ( .A(KEYINPUT91), .B(G107), .Z(n473) );
  XNOR2_X1 U464 ( .A(n472), .B(n471), .ZN(n474) );
  INV_X1 U465 ( .A(G101), .ZN(n471) );
  XNOR2_X1 U466 ( .A(n466), .B(G122), .ZN(n446) );
  XOR2_X1 U467 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n466) );
  XNOR2_X1 U468 ( .A(G128), .B(KEYINPUT24), .ZN(n516) );
  XNOR2_X1 U469 ( .A(G116), .B(G134), .ZN(n484) );
  XOR2_X1 U470 ( .A(G122), .B(G107), .Z(n485) );
  XNOR2_X1 U471 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n486) );
  XOR2_X1 U472 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n487) );
  XOR2_X1 U473 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n491) );
  XNOR2_X1 U474 ( .A(n504), .B(n385), .ZN(n682) );
  XNOR2_X1 U475 ( .A(n502), .B(n386), .ZN(n385) );
  XNOR2_X1 U476 ( .A(n503), .B(n387), .ZN(n386) );
  INV_X1 U477 ( .A(KEYINPUT70), .ZN(n412) );
  NOR2_X1 U478 ( .A1(n579), .A2(n637), .ZN(n391) );
  XNOR2_X1 U479 ( .A(n605), .B(n604), .ZN(n620) );
  NOR2_X1 U480 ( .A1(n646), .A2(n628), .ZN(n629) );
  XNOR2_X1 U481 ( .A(n647), .B(n558), .ZN(n656) );
  INV_X1 U482 ( .A(KEYINPUT6), .ZN(n558) );
  XOR2_X1 U483 ( .A(n535), .B(n536), .Z(n694) );
  XNOR2_X1 U484 ( .A(n541), .B(n534), .ZN(n536) );
  XNOR2_X1 U485 ( .A(n675), .B(KEYINPUT80), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n613), .B(KEYINPUT85), .ZN(n614) );
  XNOR2_X1 U487 ( .A(n400), .B(KEYINPUT32), .ZN(n758) );
  NAND2_X1 U488 ( .A1(n398), .A2(n365), .ZN(n396) );
  XNOR2_X1 U489 ( .A(n552), .B(KEYINPUT104), .ZN(n712) );
  BUF_X1 U490 ( .A(n698), .Z(n405) );
  XNOR2_X1 U491 ( .A(n732), .B(n733), .ZN(n402) );
  INV_X1 U492 ( .A(KEYINPUT60), .ZN(n409) );
  XNOR2_X1 U493 ( .A(n448), .B(n447), .ZN(n726) );
  XNOR2_X1 U494 ( .A(n725), .B(n724), .ZN(n447) );
  INV_X1 U495 ( .A(KEYINPUT56), .ZN(n449) );
  XNOR2_X1 U496 ( .A(n677), .B(n406), .ZN(G75) );
  INV_X1 U497 ( .A(KEYINPUT53), .ZN(n406) );
  NAND2_X1 U498 ( .A1(n430), .A2(n429), .ZN(n677) );
  NOR2_X1 U499 ( .A1(n676), .A2(G953), .ZN(n429) );
  INV_X1 U500 ( .A(n439), .ZN(n722) );
  XOR2_X1 U501 ( .A(n517), .B(n516), .Z(n360) );
  XNOR2_X1 U502 ( .A(G137), .B(G140), .ZN(n361) );
  XOR2_X1 U503 ( .A(KEYINPUT77), .B(n635), .Z(n362) );
  AND2_X1 U504 ( .A1(n439), .A2(n721), .ZN(n363) );
  XOR2_X1 U505 ( .A(n476), .B(n456), .Z(n364) );
  AND2_X1 U506 ( .A1(n397), .A2(n639), .ZN(n365) );
  NOR2_X1 U507 ( .A1(n682), .A2(G902), .ZN(n366) );
  XOR2_X1 U508 ( .A(n694), .B(n693), .Z(n367) );
  XOR2_X1 U509 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n368) );
  AND2_X1 U510 ( .A1(n371), .A2(n369), .ZN(n643) );
  NAND2_X1 U511 ( .A1(n370), .A2(KEYINPUT44), .ZN(n662) );
  NAND2_X1 U512 ( .A1(n370), .A2(n631), .ZN(n640) );
  INV_X1 U513 ( .A(n371), .ZN(n370) );
  XNOR2_X1 U514 ( .A(n371), .B(G122), .ZN(G24) );
  XNOR2_X2 U515 ( .A(n452), .B(n368), .ZN(n371) );
  XNOR2_X2 U516 ( .A(n375), .B(n664), .ZN(n392) );
  NAND2_X1 U517 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X2 U518 ( .A1(n379), .A2(n415), .ZN(n377) );
  XNOR2_X1 U519 ( .A(n380), .B(KEYINPUT18), .ZN(n421) );
  NAND2_X1 U520 ( .A1(n526), .A2(G214), .ZN(n500) );
  INV_X1 U521 ( .A(n580), .ZN(n384) );
  INV_X1 U522 ( .A(n596), .ZN(n388) );
  NAND2_X1 U523 ( .A1(n665), .A2(n392), .ZN(n667) );
  NAND2_X1 U524 ( .A1(n674), .A2(n392), .ZN(n679) );
  NAND2_X1 U525 ( .A1(n392), .A2(n753), .ZN(n735) );
  XNOR2_X1 U526 ( .A(n393), .B(n441), .ZN(n440) );
  NAND2_X1 U527 ( .A1(n394), .A2(n399), .ZN(n398) );
  INV_X1 U528 ( .A(n655), .ZN(n394) );
  NAND2_X1 U529 ( .A1(n362), .A2(n636), .ZN(n401) );
  AND2_X1 U530 ( .A1(n655), .A2(KEYINPUT106), .ZN(n395) );
  NAND2_X1 U531 ( .A1(n637), .A2(KEYINPUT106), .ZN(n397) );
  NOR2_X1 U532 ( .A1(n655), .A2(n401), .ZN(n400) );
  XNOR2_X2 U533 ( .A(n414), .B(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U534 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X2 U535 ( .A(n404), .B(n403), .ZN(n655) );
  NAND2_X1 U536 ( .A1(n642), .A2(n643), .ZN(n644) );
  NOR2_X1 U537 ( .A1(n402), .A2(n734), .ZN(G66) );
  NAND2_X1 U538 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n629), .B(KEYINPUT34), .ZN(n453) );
  NOR2_X2 U540 ( .A1(n649), .A2(n419), .ZN(n404) );
  NOR2_X2 U541 ( .A1(n546), .A2(n588), .ZN(n557) );
  NAND2_X1 U542 ( .A1(n453), .A2(n630), .ZN(n452) );
  XNOR2_X1 U543 ( .A(n442), .B(KEYINPUT96), .ZN(n648) );
  NAND2_X1 U544 ( .A1(n457), .A2(n407), .ZN(n525) );
  NAND2_X1 U545 ( .A1(n408), .A2(n364), .ZN(n407) );
  INV_X1 U546 ( .A(n495), .ZN(n408) );
  XNOR2_X1 U547 ( .A(n410), .B(n409), .ZN(G60) );
  NAND2_X1 U548 ( .A1(n688), .A2(n723), .ZN(n410) );
  XNOR2_X1 U549 ( .A(n411), .B(n367), .ZN(n461) );
  NAND2_X1 U550 ( .A1(n416), .A2(n680), .ZN(n411) );
  NAND2_X1 U551 ( .A1(n413), .A2(n680), .ZN(n686) );
  NAND2_X1 U552 ( .A1(n644), .A2(n663), .ZN(n415) );
  AND2_X1 U553 ( .A1(n681), .A2(G472), .ZN(n416) );
  NAND2_X1 U554 ( .A1(n417), .A2(n680), .ZN(n692) );
  AND2_X1 U555 ( .A1(n681), .A2(G210), .ZN(n417) );
  NAND2_X1 U556 ( .A1(n418), .A2(G217), .ZN(n732) );
  NAND2_X1 U557 ( .A1(n418), .A2(G478), .ZN(n728) );
  NAND2_X1 U558 ( .A1(n418), .A2(G469), .ZN(n448) );
  XNOR2_X2 U559 ( .A(n627), .B(KEYINPUT0), .ZN(n649) );
  XNOR2_X1 U560 ( .A(n422), .B(KEYINPUT46), .ZN(n617) );
  NAND2_X1 U561 ( .A1(n620), .A2(n712), .ZN(n423) );
  NOR2_X1 U562 ( .A1(n592), .A2(n424), .ZN(n425) );
  NAND2_X1 U563 ( .A1(n359), .A2(n593), .ZN(n424) );
  NAND2_X1 U564 ( .A1(n426), .A2(n425), .ZN(n604) );
  INV_X1 U565 ( .A(n645), .ZN(n426) );
  NOR2_X1 U566 ( .A1(n592), .A2(n428), .ZN(n427) );
  NAND2_X1 U567 ( .A1(n426), .A2(n427), .ZN(n602) );
  INV_X1 U568 ( .A(n593), .ZN(n428) );
  NAND2_X1 U569 ( .A1(n618), .A2(n438), .ZN(n437) );
  INV_X1 U570 ( .A(KEYINPUT48), .ZN(n438) );
  XNOR2_X1 U571 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U572 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U573 ( .A(n470), .B(n740), .ZN(n479) );
  NAND2_X1 U574 ( .A1(n445), .A2(n654), .ZN(n444) );
  XNOR2_X1 U575 ( .A(n653), .B(KEYINPUT99), .ZN(n445) );
  XNOR2_X1 U576 ( .A(n450), .B(n449), .ZN(G51) );
  NAND2_X1 U577 ( .A1(n451), .A2(n723), .ZN(n450) );
  XNOR2_X1 U578 ( .A(n692), .B(n691), .ZN(n451) );
  XNOR2_X2 U579 ( .A(n455), .B(n454), .ZN(n587) );
  XNOR2_X2 U580 ( .A(n475), .B(G143), .ZN(n495) );
  NOR2_X1 U581 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U582 ( .A(KEYINPUT19), .B(KEYINPUT67), .Z(n459) );
  AND2_X1 U583 ( .A1(G227), .A2(n753), .ZN(n460) );
  XNOR2_X1 U584 ( .A(n463), .B(n462), .ZN(n465) );
  INV_X1 U585 ( .A(n525), .ZN(n477) );
  XNOR2_X1 U586 ( .A(n747), .B(n361), .ZN(n514) );
  INV_X1 U587 ( .A(KEYINPUT36), .ZN(n613) );
  XNOR2_X1 U588 ( .A(n479), .B(n478), .ZN(n689) );
  INV_X1 U589 ( .A(G472), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U591 ( .A(KEYINPUT40), .ZN(n606) );
  NOR2_X1 U592 ( .A1(n648), .A2(n647), .ZN(n698) );
  INV_X1 U593 ( .A(KEYINPUT3), .ZN(n462) );
  XOR2_X1 U594 ( .A(KEYINPUT69), .B(G119), .Z(n464) );
  NAND2_X1 U595 ( .A1(G224), .A2(n753), .ZN(n468) );
  XNOR2_X2 U596 ( .A(G128), .B(KEYINPUT66), .ZN(n475) );
  XNOR2_X1 U597 ( .A(n480), .B(KEYINPUT90), .ZN(n509) );
  INV_X1 U598 ( .A(n509), .ZN(n678) );
  NAND2_X1 U599 ( .A1(G210), .A2(n483), .ZN(n481) );
  XNOR2_X2 U600 ( .A(n482), .B(n481), .ZN(n596) );
  XOR2_X1 U601 ( .A(n596), .B(KEYINPUT38), .Z(n603) );
  NAND2_X1 U602 ( .A1(G214), .A2(n483), .ZN(n590) );
  NAND2_X1 U603 ( .A1(n359), .A2(n590), .ZN(n554) );
  XNOR2_X1 U604 ( .A(n485), .B(n484), .ZN(n489) );
  XNOR2_X1 U605 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U606 ( .A(n489), .B(n488), .Z(n493) );
  NAND2_X1 U607 ( .A1(G234), .A2(n753), .ZN(n490) );
  XNOR2_X1 U608 ( .A(n491), .B(n490), .ZN(n515) );
  NAND2_X1 U609 ( .A1(G217), .A2(n515), .ZN(n492) );
  XNOR2_X1 U610 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U611 ( .A(n495), .B(n494), .ZN(n727) );
  NOR2_X1 U612 ( .A1(G902), .A2(n727), .ZN(n496) );
  XOR2_X1 U613 ( .A(G478), .B(n496), .Z(n553) );
  INV_X1 U614 ( .A(n553), .ZN(n595) );
  XNOR2_X1 U615 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n505) );
  XNOR2_X1 U616 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U617 ( .A(n747), .B(n499), .ZN(n504) );
  XNOR2_X1 U618 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U619 ( .A(n505), .B(n366), .ZN(n506) );
  XNOR2_X1 U620 ( .A(G475), .B(n506), .ZN(n594) );
  NAND2_X1 U621 ( .A1(n595), .A2(n594), .ZN(n632) );
  NOR2_X1 U622 ( .A1(n554), .A2(n632), .ZN(n508) );
  XNOR2_X1 U623 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n507) );
  XNOR2_X1 U624 ( .A(n508), .B(n507), .ZN(n608) );
  INV_X1 U625 ( .A(n608), .ZN(n570) );
  XNOR2_X1 U626 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n549) );
  XOR2_X1 U627 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n523) );
  XOR2_X1 U628 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n512) );
  NAND2_X1 U629 ( .A1(n509), .A2(G234), .ZN(n510) );
  XNOR2_X1 U630 ( .A(KEYINPUT20), .B(n510), .ZN(n520) );
  NAND2_X1 U631 ( .A1(n520), .A2(G217), .ZN(n511) );
  XNOR2_X1 U632 ( .A(n512), .B(n511), .ZN(n519) );
  NAND2_X1 U633 ( .A1(G221), .A2(n515), .ZN(n518) );
  XOR2_X1 U634 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n517) );
  NAND2_X1 U635 ( .A1(G221), .A2(n520), .ZN(n521) );
  XNOR2_X1 U636 ( .A(n521), .B(KEYINPUT21), .ZN(n633) );
  NAND2_X1 U637 ( .A1(n659), .A2(n633), .ZN(n522) );
  XNOR2_X1 U638 ( .A(n523), .B(n522), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n526), .A2(G210), .ZN(n527) );
  XNOR2_X1 U640 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U641 ( .A(n529), .B(G101), .Z(n533) );
  XNOR2_X1 U642 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X2 U643 ( .A(n538), .B(n537), .ZN(n647) );
  INV_X1 U644 ( .A(n647), .ZN(n638) );
  NAND2_X1 U645 ( .A1(n539), .A2(n638), .ZN(n540) );
  XNOR2_X1 U646 ( .A(n540), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U647 ( .A(n587), .B(KEYINPUT1), .ZN(n546) );
  BUF_X1 U648 ( .A(n546), .Z(n661) );
  NAND2_X1 U649 ( .A1(n661), .A2(n588), .ZN(n543) );
  XNOR2_X1 U650 ( .A(KEYINPUT50), .B(n543), .ZN(n544) );
  NAND2_X1 U651 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U652 ( .A1(n647), .A2(n557), .ZN(n650) );
  NAND2_X1 U653 ( .A1(n547), .A2(n650), .ZN(n548) );
  XNOR2_X1 U654 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U655 ( .A1(n570), .A2(n550), .ZN(n563) );
  NOR2_X1 U656 ( .A1(n359), .A2(n590), .ZN(n551) );
  NOR2_X1 U657 ( .A1(n632), .A2(n551), .ZN(n556) );
  NOR2_X1 U658 ( .A1(n594), .A2(n553), .ZN(n552) );
  AND2_X1 U659 ( .A1(n553), .A2(n594), .ZN(n714) );
  NOR2_X1 U660 ( .A1(n712), .A2(n714), .ZN(n583) );
  NOR2_X1 U661 ( .A1(n583), .A2(n554), .ZN(n555) );
  NOR2_X1 U662 ( .A1(n556), .A2(n555), .ZN(n561) );
  XNOR2_X1 U663 ( .A(n557), .B(KEYINPUT107), .ZN(n559) );
  INV_X1 U664 ( .A(n656), .ZN(n635) );
  XNOR2_X1 U665 ( .A(KEYINPUT33), .B(n560), .ZN(n628) );
  BUF_X1 U666 ( .A(n628), .Z(n571) );
  NOR2_X1 U667 ( .A1(n561), .A2(n571), .ZN(n562) );
  NOR2_X1 U668 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U669 ( .A(KEYINPUT119), .B(n564), .ZN(n565) );
  XNOR2_X1 U670 ( .A(n565), .B(KEYINPUT52), .ZN(n568) );
  XNOR2_X1 U671 ( .A(n566), .B(KEYINPUT14), .ZN(n575) );
  NAND2_X1 U672 ( .A1(G952), .A2(n575), .ZN(n567) );
  XOR2_X1 U673 ( .A(KEYINPUT92), .B(n567), .Z(n574) );
  NAND2_X1 U674 ( .A1(n568), .A2(n574), .ZN(n569) );
  XNOR2_X1 U675 ( .A(n569), .B(KEYINPUT120), .ZN(n573) );
  OR2_X1 U676 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U677 ( .A1(n573), .A2(n572), .ZN(n676) );
  INV_X1 U678 ( .A(KEYINPUT78), .ZN(n668) );
  INV_X1 U679 ( .A(n661), .ZN(n637) );
  NAND2_X1 U680 ( .A1(n753), .A2(n574), .ZN(n624) );
  NAND2_X1 U681 ( .A1(G902), .A2(n575), .ZN(n621) );
  NOR2_X1 U682 ( .A1(G900), .A2(n621), .ZN(n576) );
  NAND2_X1 U683 ( .A1(G953), .A2(n576), .ZN(n577) );
  NAND2_X1 U684 ( .A1(n624), .A2(n577), .ZN(n593) );
  NAND2_X1 U685 ( .A1(n659), .A2(n593), .ZN(n578) );
  NOR2_X1 U686 ( .A1(n633), .A2(n578), .ZN(n580) );
  NAND2_X1 U687 ( .A1(n590), .A2(n610), .ZN(n579) );
  INV_X1 U688 ( .A(KEYINPUT72), .ZN(n586) );
  NOR2_X1 U689 ( .A1(n586), .A2(KEYINPUT47), .ZN(n585) );
  AND2_X1 U690 ( .A1(n647), .A2(n580), .ZN(n581) );
  XOR2_X1 U691 ( .A(KEYINPUT28), .B(n581), .Z(n582) );
  NOR2_X1 U692 ( .A1(n582), .A2(n587), .ZN(n607) );
  AND2_X1 U693 ( .A1(n626), .A2(n607), .ZN(n709) );
  INV_X1 U694 ( .A(n583), .ZN(n654) );
  NAND2_X1 U695 ( .A1(n709), .A2(n654), .ZN(n584) );
  XNOR2_X1 U696 ( .A(n585), .B(n584), .ZN(n601) );
  NAND2_X1 U697 ( .A1(n586), .A2(KEYINPUT47), .ZN(n599) );
  XNOR2_X1 U698 ( .A(n589), .B(KEYINPUT95), .ZN(n645) );
  NAND2_X1 U699 ( .A1(n647), .A2(n590), .ZN(n591) );
  XNOR2_X1 U700 ( .A(KEYINPUT30), .B(n591), .ZN(n592) );
  NOR2_X1 U701 ( .A1(n595), .A2(n594), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n596), .A2(n630), .ZN(n597) );
  NOR2_X1 U703 ( .A1(n602), .A2(n597), .ZN(n707) );
  XNOR2_X1 U704 ( .A(KEYINPUT79), .B(n707), .ZN(n598) );
  AND2_X1 U705 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U706 ( .A1(n601), .A2(n600), .ZN(n619) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(KEYINPUT39), .Z(n605) );
  XOR2_X1 U708 ( .A(KEYINPUT42), .B(n609), .Z(n759) );
  INV_X1 U709 ( .A(n610), .ZN(n612) );
  NOR2_X1 U710 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U711 ( .A1(n637), .A2(n616), .ZN(n718) );
  NAND2_X1 U712 ( .A1(n617), .A2(n718), .ZN(n618) );
  NAND2_X1 U713 ( .A1(n714), .A2(n620), .ZN(n721) );
  NOR2_X1 U714 ( .A1(n668), .A2(n751), .ZN(n665) );
  INV_X1 U715 ( .A(n621), .ZN(n622) );
  NOR2_X1 U716 ( .A1(G898), .A2(n753), .ZN(n743) );
  NAND2_X1 U717 ( .A1(n622), .A2(n743), .ZN(n623) );
  NAND2_X1 U718 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U719 ( .A(KEYINPUT83), .ZN(n631) );
  INV_X1 U720 ( .A(n632), .ZN(n634) );
  AND2_X1 U721 ( .A1(n637), .A2(n659), .ZN(n636) );
  AND2_X1 U722 ( .A1(n659), .A2(n638), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n642), .ZN(n641) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n652) );
  XOR2_X1 U725 ( .A(KEYINPUT31), .B(KEYINPUT98), .Z(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n715) );
  NOR2_X1 U727 ( .A1(n698), .A2(n715), .ZN(n653) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U729 ( .A(KEYINPUT82), .B(n657), .Z(n658) );
  NOR2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n696) );
  NAND2_X1 U732 ( .A1(n662), .A2(KEYINPUT83), .ZN(n663) );
  XNOR2_X1 U733 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n664) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n666) );
  NAND2_X2 U735 ( .A1(n667), .A2(n666), .ZN(n681) );
  NAND2_X1 U736 ( .A1(n668), .A2(n721), .ZN(n671) );
  NAND2_X1 U737 ( .A1(n721), .A2(KEYINPUT2), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n669), .A2(KEYINPUT78), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U741 ( .A1(n681), .A2(n679), .ZN(n675) );
  AND2_X2 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n684) );
  XNOR2_X1 U744 ( .A(n682), .B(KEYINPUT88), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U746 ( .A(n686), .B(n685), .ZN(n688) );
  NOR2_X1 U747 ( .A1(G952), .A2(n753), .ZN(n687) );
  XNOR2_X1 U748 ( .A(KEYINPUT89), .B(n687), .ZN(n723) );
  XNOR2_X1 U749 ( .A(n689), .B(KEYINPUT55), .ZN(n690) );
  XOR2_X1 U750 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n693) );
  NAND2_X1 U751 ( .A1(n461), .A2(n723), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n695), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U753 ( .A(G101), .B(n696), .ZN(G3) );
  NAND2_X1 U754 ( .A1(n712), .A2(n405), .ZN(n697) );
  XNOR2_X1 U755 ( .A(n697), .B(G104), .ZN(G6) );
  XNOR2_X1 U756 ( .A(G107), .B(KEYINPUT110), .ZN(n702) );
  XOR2_X1 U757 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n700) );
  NAND2_X1 U758 ( .A1(n405), .A2(n714), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U760 ( .A(n702), .B(n701), .ZN(G9) );
  XOR2_X1 U761 ( .A(G110), .B(n703), .Z(G12) );
  XOR2_X1 U762 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n705) );
  NAND2_X1 U763 ( .A1(n709), .A2(n714), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U765 ( .A(G128), .B(n706), .Z(G30) );
  XOR2_X1 U766 ( .A(G143), .B(n707), .Z(n708) );
  XNOR2_X1 U767 ( .A(KEYINPUT112), .B(n708), .ZN(G45) );
  XOR2_X1 U768 ( .A(G146), .B(KEYINPUT113), .Z(n711) );
  NAND2_X1 U769 ( .A1(n709), .A2(n712), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(G48) );
  NAND2_X1 U771 ( .A1(n715), .A2(n712), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n713), .B(G113), .ZN(G15) );
  NAND2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U774 ( .A(n716), .B(G116), .ZN(G18) );
  XOR2_X1 U775 ( .A(KEYINPUT114), .B(KEYINPUT37), .Z(n717) );
  XNOR2_X1 U776 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U777 ( .A(G125), .B(n719), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(KEYINPUT115), .Z(n720) );
  XNOR2_X1 U779 ( .A(n721), .B(n720), .ZN(G36) );
  XOR2_X1 U780 ( .A(G140), .B(n722), .Z(G42) );
  INV_X1 U781 ( .A(n723), .ZN(n734) );
  XOR2_X1 U782 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  NOR2_X1 U783 ( .A1(n734), .A2(n726), .ZN(G54) );
  XNOR2_X1 U784 ( .A(n727), .B(KEYINPUT122), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n734), .A2(n730), .ZN(G63) );
  XOR2_X1 U787 ( .A(n731), .B(KEYINPUT123), .Z(n733) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT124), .ZN(n739) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n746) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U795 ( .A(KEYINPUT125), .B(n744), .Z(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(n752) );
  XNOR2_X1 U798 ( .A(G227), .B(n752), .ZN(n749) );
  NAND2_X1 U799 ( .A1(G900), .A2(n749), .ZN(n750) );
  NAND2_X1 U800 ( .A1(n750), .A2(G953), .ZN(n756) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G72) );
  XOR2_X1 U804 ( .A(G119), .B(KEYINPUT126), .Z(n757) );
  XNOR2_X1 U805 ( .A(n758), .B(n757), .ZN(G21) );
  XNOR2_X1 U806 ( .A(G137), .B(KEYINPUT127), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n760), .B(n759), .ZN(G39) );
  XOR2_X1 U808 ( .A(n761), .B(G131), .Z(G33) );
endmodule

