//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n201), .B(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G223), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(new_n248), .ZN(new_n252));
  INV_X1    g0052(.A(G222), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n244), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n250), .B1(new_n251), .B2(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G274), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(KEYINPUT66), .B(G226), .Z(new_n266));
  OAI211_X1 g0066(.A(new_n259), .B(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(G200), .B2(new_n267), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n216), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n206), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(G50), .ZN(new_n278));
  INV_X1    g0078(.A(new_n275), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n207), .A2(G33), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n279), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n285), .B2(KEYINPUT67), .ZN(new_n286));
  OR2_X1    g0086(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n270), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n267), .A2(G169), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n267), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n288), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G20), .A2(G77), .ZN(new_n299));
  INV_X1    g0099(.A(new_n283), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT15), .B(G87), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n299), .B1(new_n280), .B2(new_n300), .C1(new_n281), .C2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(new_n275), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n272), .A2(new_n251), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n277), .B2(new_n251), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n249), .A2(G238), .ZN(new_n307));
  INV_X1    g0107(.A(G107), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n307), .B1(new_n308), .B2(new_n252), .C1(new_n309), .C2(new_n254), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n258), .ZN(new_n311));
  INV_X1    g0111(.A(new_n265), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n312), .A2(G244), .B1(G274), .B2(new_n262), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT68), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT68), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G200), .ZN(new_n319));
  AOI21_X1  g0119(.A(G190), .B1(new_n315), .B2(new_n317), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n306), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(G179), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(G169), .A3(new_n317), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n306), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n298), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(KEYINPUT7), .B1(new_n330), .B2(new_n207), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n248), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G68), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n337), .B2(new_n201), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n283), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n327), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n247), .A2(new_n207), .A3(new_n248), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n336), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n340), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n275), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n280), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n272), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n277), .B2(new_n349), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(G223), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n353));
  OAI211_X1 g0153(.A(G226), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n354));
  INV_X1    g0154(.A(G87), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n353), .B(new_n354), .C1(new_n246), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n258), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n263), .B1(new_n265), .B2(new_n309), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n268), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n356), .B2(new_n258), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(G200), .B2(new_n361), .ZN(new_n362));
  AND4_X1   g0162(.A1(KEYINPUT73), .A2(new_n348), .A3(new_n352), .A4(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT16), .B1(new_n346), .B2(new_n340), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n334), .A2(new_n327), .A3(new_n341), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n351), .B1(new_n366), .B2(new_n275), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT73), .B1(new_n367), .B2(new_n362), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT17), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n361), .A2(G179), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n361), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n279), .B1(new_n364), .B2(new_n365), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(new_n351), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n374), .B(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT17), .B1(new_n367), .B2(new_n362), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n257), .A2(G238), .A3(new_n264), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n263), .ZN(new_n382));
  OAI211_X1 g0182(.A(G226), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n383));
  OAI211_X1 g0183(.A(G232), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G33), .A2(G97), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT13), .B(new_n382), .C1(new_n258), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n258), .ZN(new_n389));
  INV_X1    g0189(.A(new_n382), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(G169), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT14), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n393), .A2(KEYINPUT72), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI221_X1 g0195(.A(G169), .B1(KEYINPUT72), .B2(new_n393), .C1(new_n387), .C2(new_n391), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(KEYINPUT69), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n382), .B1(new_n386), .B2(new_n258), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n388), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT69), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n398), .B2(new_n388), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n397), .A2(G179), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n396), .A3(new_n402), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n281), .A2(new_n251), .B1(new_n207), .B2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT70), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n202), .B2(new_n300), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n404), .A2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n275), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g0208(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n408), .B(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G13), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(G1), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(G20), .A3(new_n336), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT12), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n336), .B2(new_n277), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(G200), .B1(new_n387), .B2(new_n391), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n417), .B(new_n420), .C1(new_n268), .C2(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n326), .A2(new_n380), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(G238), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n426));
  OAI211_X1 g0226(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G116), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n258), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n261), .A2(G1), .ZN(new_n431));
  INV_X1    g0231(.A(G250), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G274), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n261), .A2(new_n434), .A3(G1), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n257), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n268), .ZN(new_n438));
  AOI21_X1  g0238(.A(G20), .B1(new_n247), .B2(new_n248), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G68), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT77), .B(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G20), .B2(new_n385), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n207), .B1(new_n441), .B2(new_n385), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n355), .A2(new_n446), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n445), .A2(KEYINPUT78), .B1(G107), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  INV_X1    g0249(.A(new_n385), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(KEYINPUT77), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(KEYINPUT77), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n454), .B2(new_n207), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n444), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n275), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n437), .A2(G200), .ZN(new_n458));
  INV_X1    g0258(.A(new_n301), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(new_n271), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n206), .A2(G33), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n271), .A2(new_n462), .A3(new_n216), .A4(new_n274), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G87), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n457), .A2(new_n458), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n456), .B2(new_n275), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT80), .A3(new_n458), .A4(new_n465), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n438), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n437), .A2(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n295), .B2(new_n437), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n464), .A2(new_n459), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n447), .A2(G107), .ZN(new_n476));
  XOR2_X1   g0276(.A(KEYINPUT77), .B(KEYINPUT19), .Z(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n477), .B2(new_n450), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n478), .B2(new_n449), .ZN(new_n479));
  INV_X1    g0279(.A(new_n455), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n443), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n461), .B(new_n475), .C1(new_n481), .C2(new_n279), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n469), .A2(new_n484), .A3(new_n475), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n474), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n471), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n431), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(new_n490), .A2(new_n434), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT81), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n490), .A2(new_n492), .A3(G270), .A4(new_n257), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G264), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n495));
  OAI211_X1 g0295(.A(G257), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n496));
  XOR2_X1   g0296(.A(KEYINPUT82), .B(G303), .Z(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n252), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n258), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n490), .A2(G270), .A3(new_n257), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT21), .A3(G169), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n494), .A2(G179), .A3(new_n499), .A4(new_n501), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT20), .ZN(new_n505));
  INV_X1    g0305(.A(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n207), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n446), .B2(G33), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n507), .B1(new_n509), .B2(new_n207), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n505), .B1(new_n510), .B2(new_n279), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n246), .A2(G97), .ZN(new_n512));
  AOI21_X1  g0312(.A(G20), .B1(new_n512), .B2(new_n508), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT20), .B(new_n275), .C1(new_n513), .C2(new_n507), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n271), .A2(new_n506), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n464), .B2(new_n506), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT83), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(KEYINPUT83), .A3(new_n517), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n503), .A2(new_n504), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n515), .A2(KEYINPUT83), .A3(new_n517), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n518), .ZN(new_n523));
  INV_X1    g0323(.A(G200), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n501), .A2(new_n493), .A3(new_n491), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n498), .A2(new_n258), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n494), .A2(new_n268), .A3(new_n499), .A4(new_n501), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G169), .B1(new_n525), .B2(new_n526), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n519), .B2(new_n520), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT84), .B1(new_n532), .B2(KEYINPUT21), .ZN(new_n533));
  OAI211_X1 g0333(.A(G169), .B(new_n502), .C1(new_n522), .C2(new_n518), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT84), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT21), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI211_X1 g0337(.A(new_n521), .B(new_n530), .C1(new_n533), .C2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n490), .A2(new_n257), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G257), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n491), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT75), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT4), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(KEYINPUT4), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n543), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n249), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n541), .B1(new_n550), .B2(new_n258), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n272), .A2(G97), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(G97), .B2(new_n463), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n555), .A2(new_n446), .A3(G107), .ZN(new_n556));
  XNOR2_X1  g0356(.A(G97), .B(G107), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n558), .A2(new_n207), .B1(new_n251), .B2(new_n300), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n308), .B1(new_n345), .B2(new_n332), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n275), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT74), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n275), .C1(new_n559), .C2(new_n560), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n554), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n549), .A2(new_n548), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n258), .B1(new_n566), .B2(new_n546), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n540), .A2(new_n491), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT76), .B1(new_n569), .B2(G200), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT76), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n571), .B(new_n524), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n552), .B(new_n565), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G250), .B(new_n244), .C1(new_n328), .C2(new_n329), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n575));
  INV_X1    g0375(.A(G294), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n575), .C1(new_n246), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n258), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n539), .A2(G264), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n491), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n295), .B2(new_n580), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n308), .A2(KEYINPUT23), .A3(G20), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT23), .B1(new_n308), .B2(G20), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(G20), .B2(new_n428), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n207), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n252), .A2(new_n590), .A3(new_n207), .A4(G87), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n584), .B(new_n587), .C1(new_n589), .C2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n583), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(KEYINPUT86), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n593), .B2(new_n583), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n279), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n413), .A2(G20), .A3(new_n308), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n599), .A2(KEYINPUT25), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(KEYINPUT25), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n600), .B(new_n601), .C1(new_n308), .C2(new_n463), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n582), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n562), .A2(new_n564), .ZN(new_n604));
  INV_X1    g0404(.A(new_n554), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n567), .A2(new_n568), .A3(G179), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n551), .B2(new_n371), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n580), .A2(new_n524), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT87), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n580), .A2(new_n612), .A3(new_n524), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n580), .A2(G190), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n589), .A2(new_n591), .ZN(new_n616));
  OAI211_X1 g0416(.A(KEYINPUT86), .B(new_n584), .C1(new_n616), .C2(new_n587), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n593), .A2(new_n583), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n597), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n602), .B1(new_n619), .B2(new_n275), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n573), .A2(new_n603), .A3(new_n609), .A4(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n425), .A2(new_n487), .A3(new_n538), .A4(new_n622), .ZN(G372));
  AOI22_X1  g0423(.A1(new_n325), .A2(new_n422), .B1(new_n418), .B2(new_n403), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n348), .A2(new_n352), .A3(new_n362), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT73), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n367), .A2(KEYINPUT73), .A3(new_n362), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n377), .B1(new_n629), .B2(KEYINPUT17), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n376), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n293), .B1(new_n288), .B2(new_n296), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n482), .A2(new_n473), .ZN(new_n634));
  INV_X1    g0434(.A(new_n521), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n532), .A2(KEYINPUT84), .A3(KEYINPUT21), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n603), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n634), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n466), .A2(new_n438), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n573), .A3(new_n609), .A4(new_n621), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n634), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n606), .A2(KEYINPUT88), .A3(new_n608), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT88), .B1(new_n606), .B2(new_n608), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n642), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n471), .A2(new_n486), .A3(new_n609), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n645), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n633), .B1(new_n424), .B2(new_n651), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n533), .A2(new_n537), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n413), .A2(new_n207), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT89), .Z(new_n656));
  INV_X1    g0456(.A(G213), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n654), .B2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n523), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n653), .A2(new_n635), .A3(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n664), .B(G330), .C1(new_n538), .C2(new_n663), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT90), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT90), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n621), .B1(new_n620), .B2(new_n662), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n603), .ZN(new_n671));
  INV_X1    g0471(.A(new_n603), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n662), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n661), .B1(new_n653), .B2(new_n635), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n671), .A3(new_n673), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n673), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n210), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n447), .A2(G107), .A3(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n214), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n578), .A2(new_n579), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n502), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n437), .A2(new_n295), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n551), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n691), .A4(new_n551), .ZN(new_n695));
  AOI21_X1  g0495(.A(G179), .B1(new_n430), .B2(new_n436), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n569), .A2(new_n502), .A3(new_n580), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n661), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n622), .A2(new_n538), .A3(new_n487), .A4(new_n662), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n698), .A2(new_n661), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n699), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n704), .A2(KEYINPUT91), .A3(G330), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT91), .B1(new_n704), .B2(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n573), .A2(new_n609), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n638), .A2(new_n708), .A3(new_n621), .A4(new_n642), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n649), .A2(new_n645), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT26), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n709), .A2(new_n710), .A3(new_n712), .A4(new_n634), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .A3(new_n662), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n651), .A2(new_n661), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n707), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n688), .B1(new_n718), .B2(G1), .ZN(G364));
  NOR2_X1   g0519(.A1(new_n412), .A2(G20), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G45), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n684), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n538), .A2(new_n663), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(new_n664), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n216), .B1(G20), .B2(new_n371), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n215), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n239), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n682), .A2(new_n252), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n682), .A2(new_n330), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n740), .A2(G355), .B1(new_n506), .B2(new_n682), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n733), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n207), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n295), .A2(new_n524), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT93), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G159), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT32), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n524), .A2(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n745), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n308), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n207), .A2(new_n268), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n753), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n252), .B1(new_n757), .B2(new_n355), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n744), .A2(new_n295), .A3(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(G179), .A3(new_n524), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G77), .A2(new_n759), .B1(new_n761), .B2(G58), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n295), .A2(new_n524), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(new_n756), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n202), .B2(new_n765), .ZN(new_n766));
  OR4_X1    g0566(.A1(new_n752), .A2(new_n755), .A3(new_n758), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n747), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n763), .A2(new_n743), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n769), .A2(G97), .B1(G68), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n749), .ZN(new_n775));
  OR2_X1    g0575(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(KEYINPUT95), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G329), .ZN(new_n780));
  INV_X1    g0580(.A(G283), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n754), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n757), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n759), .A2(G311), .B1(new_n783), .B2(G303), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n771), .A2(new_n785), .B1(new_n764), .B2(G326), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n252), .B1(new_n761), .B2(G322), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n782), .B(new_n788), .C1(G294), .C2(new_n769), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n774), .B1(new_n780), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n742), .B1(new_n791), .B2(new_n731), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n722), .B1(new_n730), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n669), .B1(G330), .B2(new_n724), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n794), .B2(new_n722), .ZN(G396));
  INV_X1    g0595(.A(new_n722), .ZN(new_n796));
  INV_X1    g0596(.A(new_n731), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n726), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n252), .B1(new_n202), .B2(new_n757), .C1(new_n754), .C2(new_n336), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n761), .A2(G143), .B1(new_n771), .B2(G150), .ZN(new_n800));
  INV_X1    g0600(.A(G137), .ZN(new_n801));
  INV_X1    g0601(.A(new_n759), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n801), .B2(new_n765), .C1(new_n750), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT34), .ZN(new_n804));
  INV_X1    g0604(.A(new_n769), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n335), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n799), .B(new_n806), .C1(new_n804), .C2(new_n803), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n779), .A2(G132), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n779), .A2(G311), .ZN(new_n809));
  INV_X1    g0609(.A(new_n754), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G87), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n252), .B1(new_n761), .B2(G294), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n783), .A2(G107), .B1(new_n771), .B2(G283), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n759), .A2(G116), .B1(G303), .B2(new_n764), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G97), .B2(new_n769), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n807), .A2(new_n808), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n796), .B1(G77), .B2(new_n798), .C1(new_n817), .C2(new_n797), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n306), .B(new_n661), .C1(new_n323), .C2(new_n324), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n661), .B1(new_n303), .B2(new_n305), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n321), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n325), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n818), .B1(new_n824), .B2(new_n725), .ZN(new_n825));
  INV_X1    g0625(.A(new_n707), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n715), .B(new_n824), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n796), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G384));
  INV_X1    g0631(.A(new_n558), .ZN(new_n832));
  OAI211_X1 g0632(.A(G116), .B(new_n217), .C1(new_n832), .C2(KEYINPUT35), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(KEYINPUT35), .B2(new_n832), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT36), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n214), .A2(new_n251), .A3(new_n337), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n202), .A2(G68), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n206), .B(G13), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  INV_X1    g0640(.A(new_n659), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n841), .A2(new_n372), .B1(new_n373), .B2(new_n351), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n627), .A2(new_n628), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n627), .A2(new_n845), .A3(new_n628), .A4(new_n842), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n841), .B1(new_n373), .B2(new_n351), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI221_X4 g0648(.A(new_n840), .B1(new_n844), .B2(new_n846), .C1(new_n379), .C2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n630), .B2(new_n376), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT99), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n374), .A2(new_n625), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n847), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n374), .B2(new_n625), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n363), .A2(new_n368), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n856), .A2(KEYINPUT100), .A3(new_n845), .A4(new_n842), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT100), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n846), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n850), .B1(new_n860), .B2(KEYINPUT101), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT101), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n855), .A2(new_n857), .A3(new_n862), .A4(new_n859), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT102), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n849), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n860), .A2(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n379), .A2(new_n848), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n863), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n840), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n418), .A2(new_n661), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n419), .A2(new_n873), .A3(new_n422), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n403), .A2(new_n418), .A3(new_n661), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT97), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT97), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n403), .A2(new_n418), .A3(new_n877), .A4(new_n661), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT98), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT98), .A4(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n704), .A2(new_n883), .A3(new_n823), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n844), .A2(new_n846), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n868), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n849), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT103), .B(new_n885), .C1(new_n884), .C2(new_n889), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n872), .A2(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n425), .A2(new_n704), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n894), .B(new_n895), .Z(new_n896));
  INV_X1    g0696(.A(G330), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n889), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n662), .B(new_n823), .C1(new_n644), .C2(new_n650), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT96), .ZN(new_n901));
  INV_X1    g0701(.A(new_n819), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n899), .B(new_n883), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n376), .A2(new_n841), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n419), .A2(new_n661), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n866), .A2(new_n910), .A3(new_n871), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n899), .A2(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n633), .B1(new_n424), .B2(new_n716), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n898), .A2(new_n916), .B1(new_n206), .B2(new_n720), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n898), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n839), .B1(new_n917), .B2(new_n918), .ZN(G367));
  OAI211_X1 g0719(.A(new_n573), .B(new_n609), .C1(new_n565), .C2(new_n662), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n606), .A2(new_n608), .A3(new_n661), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT104), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(new_n678), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n609), .B1(new_n924), .B2(new_n603), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n662), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n662), .B1(new_n469), .B2(new_n465), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n634), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n642), .B2(new_n929), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n926), .A2(new_n928), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n924), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n933), .A2(new_n935), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n936), .A2(new_n675), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n936), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n676), .B2(new_n924), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n683), .B(KEYINPUT41), .Z(new_n942));
  INV_X1    g0742(.A(new_n678), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n669), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n677), .B1(new_n671), .B2(new_n673), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT106), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n943), .B1(new_n666), .B2(new_n667), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n944), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n668), .A2(new_n678), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n946), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT107), .B1(new_n953), .B2(new_n717), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT44), .B1(new_n937), .B2(new_n680), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n924), .A2(new_n956), .A3(new_n679), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n937), .A2(KEYINPUT45), .A3(new_n680), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT45), .B1(new_n937), .B2(new_n680), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n955), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT105), .B1(new_n960), .B2(new_n675), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n675), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT107), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n718), .A2(new_n964), .A3(new_n952), .A4(new_n950), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n960), .A2(KEYINPUT105), .A3(new_n675), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n954), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n942), .B1(new_n967), .B2(new_n718), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n721), .A2(G1), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n939), .B(new_n941), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n737), .A2(new_n235), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n732), .B1(new_n210), .B2(new_n301), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n754), .A2(new_n446), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n759), .A2(G283), .B1(G311), .B2(new_n764), .ZN(new_n974));
  INV_X1    g0774(.A(new_n497), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n252), .B1(new_n761), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n976), .C1(new_n749), .C2(new_n977), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n973), .B(new_n978), .C1(G107), .C2(new_n769), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n757), .B2(new_n506), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n576), .C2(new_n770), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT108), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT109), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n769), .A2(G68), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n761), .A2(G150), .B1(new_n764), .B2(G143), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT110), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n754), .A2(new_n251), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n252), .B1(new_n750), .B2(new_n770), .C1(new_n802), .C2(new_n202), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n749), .A2(new_n801), .B1(new_n335), .B2(new_n757), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(KEYINPUT111), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n994), .C1(KEYINPUT111), .C2(new_n993), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n986), .A2(KEYINPUT47), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n731), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT47), .B1(new_n986), .B2(new_n995), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n796), .B1(new_n971), .B2(new_n972), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT112), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(new_n1000), .B1(new_n727), .B2(new_n931), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n970), .A2(new_n1002), .ZN(G387));
  NAND2_X1  g0803(.A1(new_n954), .A2(new_n965), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n684), .B1(new_n953), .B2(new_n717), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n685), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n740), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(G107), .B2(new_n210), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n232), .A2(new_n261), .ZN(new_n1010));
  AOI211_X1 g0810(.A(G45), .B(new_n1007), .C1(G68), .C2(G77), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n280), .A2(G50), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n737), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1009), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n330), .B1(new_n754), .B2(new_n506), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n759), .A2(new_n975), .B1(G322), .B2(new_n764), .ZN(new_n1017));
  INV_X1    g0817(.A(G311), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n770), .C1(new_n977), .C2(new_n760), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT48), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n781), .B2(new_n805), .C1(new_n576), .C2(new_n757), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT49), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1016), .B(new_n1023), .C1(G326), .C2(new_n775), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n769), .A2(new_n459), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n202), .B2(new_n760), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT113), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n783), .A2(G77), .B1(new_n764), .B2(G159), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n330), .B1(new_n771), .B2(new_n349), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n336), .C2(new_n802), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n973), .B(new_n1031), .C1(G150), .C2(new_n775), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1024), .A2(new_n1025), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n796), .B1(new_n733), .B2(new_n1015), .C1(new_n1033), .C2(new_n797), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n674), .B2(new_n727), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT114), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n969), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1006), .B(new_n1036), .C1(new_n953), .C2(new_n1037), .ZN(G393));
  INV_X1    g0838(.A(new_n962), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n960), .A2(new_n675), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n969), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n732), .B1(new_n446), .B2(new_n210), .C1(new_n737), .C2(new_n242), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(new_n796), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n330), .B1(new_n759), .B2(new_n349), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n783), .A2(G68), .B1(new_n771), .B2(G50), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n811), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n775), .A2(G143), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n769), .A2(G77), .ZN(new_n1048));
  INV_X1    g0848(.A(G150), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n765), .A2(new_n1049), .B1(new_n760), .B2(new_n750), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT51), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n775), .A2(G322), .B1(G283), .B2(new_n783), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n330), .B1(new_n802), .B2(new_n576), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n765), .A2(new_n977), .B1(new_n760), .B2(new_n1018), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  OR4_X1    g0857(.A1(new_n755), .A2(new_n1054), .A3(new_n1055), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n769), .A2(G116), .B1(new_n975), .B2(new_n771), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT116), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1052), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n731), .B1(new_n1061), .B2(KEYINPUT117), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1043), .B1(new_n1062), .B2(new_n1063), .C1(new_n937), .C2(new_n728), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1041), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n967), .A2(new_n683), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1004), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G390));
  OAI21_X1  g0870(.A(new_n796), .B1(new_n349), .B2(new_n798), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n913), .A2(new_n726), .ZN(new_n1072));
  OAI21_X1  g0872(.A(KEYINPUT53), .B1(new_n757), .B2(new_n1049), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(KEYINPUT54), .B(G143), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n252), .C1(new_n802), .C2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n757), .A2(KEYINPUT53), .A3(new_n1049), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n810), .A2(G50), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n761), .A2(G132), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n771), .A2(G137), .B1(new_n764), .B2(G128), .ZN(new_n1080));
  AND4_X1   g0880(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(G125), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1081), .B1(new_n750), .B2(new_n805), .C1(new_n1082), .C2(new_n778), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n778), .A2(new_n576), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n765), .A2(new_n781), .B1(new_n760), .B2(new_n506), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n802), .A2(new_n446), .B1(new_n308), .B2(new_n770), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G68), .C2(new_n810), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n330), .B1(new_n757), .B2(new_n355), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT122), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n1048), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1071), .B(new_n1072), .C1(new_n731), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n821), .A2(new_n822), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n713), .A2(new_n662), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n902), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n909), .B1(new_n1095), .B2(new_n883), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n872), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n900), .A2(new_n902), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT96), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n903), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n909), .B1(new_n1100), .B2(new_n883), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1097), .B1(new_n913), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n704), .A2(G330), .A3(new_n823), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n883), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1104), .B1(new_n1099), .B2(new_n903), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n911), .B(new_n912), .C1(new_n1107), .C2(new_n909), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n823), .B(new_n883), .C1(new_n705), .C2(new_n706), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1097), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT121), .B1(new_n1111), .B2(new_n1037), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1108), .A2(new_n1097), .A3(new_n1109), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1105), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1108), .B2(new_n1097), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT121), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n969), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1092), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n904), .A2(new_n905), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n823), .B1(new_n705), .B2(new_n706), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1104), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n1114), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1103), .A2(KEYINPUT118), .A3(new_n1104), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT118), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n1095), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT119), .B1(new_n1128), .B2(new_n1109), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1095), .ZN(new_n1130));
  AND4_X1   g0930(.A1(KEYINPUT119), .A2(new_n1130), .A3(new_n1109), .A4(new_n1125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1124), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n633), .B1(new_n424), .B2(new_n716), .C1(new_n895), .C2(new_n897), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(KEYINPUT120), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT119), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT118), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1095), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1125), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1109), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1137), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1130), .A2(new_n1109), .A3(KEYINPUT119), .A4(new_n1125), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1123), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1136), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1135), .A2(new_n1147), .A3(new_n1111), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1133), .B1(new_n1149), .B2(new_n1124), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n684), .B1(new_n1116), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1119), .A2(new_n1152), .ZN(G378));
  OAI21_X1  g0953(.A(new_n796), .B1(G50), .B2(new_n798), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n289), .A2(new_n659), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n298), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n293), .B2(new_n297), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1159));
  OR3_X1    g0959(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1162), .A2(new_n726), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n330), .B2(new_n260), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n252), .C1(new_n783), .C2(G77), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n761), .A2(G107), .B1(new_n764), .B2(G116), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n759), .A2(new_n459), .B1(new_n771), .B2(G97), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n987), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n810), .A2(G58), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT123), .Z(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(G283), .C2(new_n779), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1165), .B1(new_n1173), .B2(KEYINPUT58), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n757), .A2(new_n1074), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT124), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n761), .A2(G128), .B1(new_n771), .B2(G132), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n801), .C2(new_n802), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n769), .A2(G150), .B1(G125), .B2(new_n764), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT125), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT59), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n775), .A2(G124), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n810), .C2(G159), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1174), .B1(KEYINPUT58), .B2(new_n1173), .C1(new_n1184), .C2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1154), .B(new_n1163), .C1(new_n731), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n913), .A2(new_n909), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n907), .A3(new_n906), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1162), .B1(new_n894), .B2(G330), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n892), .A2(new_n893), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n849), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n870), .B2(KEYINPUT102), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n864), .A2(new_n865), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n886), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1197), .A3(G330), .A4(new_n1162), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1192), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1193), .A2(new_n1197), .A3(G330), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1162), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n914), .A3(new_n1198), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1189), .B1(new_n1205), .B2(new_n969), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1203), .A2(new_n914), .A3(new_n1198), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n914), .B1(new_n1203), .B2(new_n1198), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1133), .B1(new_n1116), .B2(new_n1150), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n683), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1134), .B1(new_n1111), .B2(new_n1146), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1212), .B2(new_n1205), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1211), .B2(new_n1213), .ZN(G375));
  OAI21_X1  g1014(.A(new_n796), .B1(G68), .B2(new_n798), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n779), .A2(G128), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n769), .A2(G50), .ZN(new_n1217));
  INV_X1    g1017(.A(G132), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n802), .A2(new_n1049), .B1(new_n1218), .B2(new_n765), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n252), .B1(new_n760), .B2(new_n801), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n750), .A2(new_n757), .B1(new_n770), .B2(new_n1074), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1216), .A2(new_n1171), .A3(new_n1217), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1026), .B1(new_n781), .B2(new_n760), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT126), .Z(new_n1225));
  AOI22_X1  g1025(.A1(new_n759), .A2(G107), .B1(new_n771), .B2(G116), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n446), .B2(new_n757), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n330), .B1(new_n765), .B2(new_n576), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1227), .A2(new_n991), .A3(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G303), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n778), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1223), .B1(new_n1225), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1215), .B1(new_n1232), .B2(new_n731), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n883), .B2(new_n726), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1146), .B2(new_n1037), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT127), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT127), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n1234), .C1(new_n1146), .C2(new_n1037), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n942), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1149), .A2(new_n1133), .A3(new_n1124), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1135), .A2(new_n1147), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n970), .A2(new_n1069), .A3(new_n1002), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G393), .A2(G396), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1244), .A2(new_n1245), .A3(G381), .A4(G384), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(G407));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1246), .B2(new_n660), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(G213), .ZN(G409));
  XOR2_X1   g1050(.A(G393), .B(G396), .Z(new_n1251));
  AND3_X1   g1051(.A1(new_n970), .A2(new_n1002), .A3(new_n1069), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1069), .B1(new_n970), .B2(new_n1002), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(G390), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(G396), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1244), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1212), .A2(new_n1240), .A3(new_n1205), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1206), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1152), .A3(new_n1119), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1119), .A2(new_n1152), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(G375), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1150), .A2(new_n684), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1241), .A2(KEYINPUT60), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1265), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1269), .A2(new_n1239), .A3(G384), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G384), .B1(new_n1269), .B2(new_n1239), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n657), .A2(G343), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1263), .A2(new_n1264), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G378), .B(new_n1206), .C1(new_n1213), .C2(new_n1211), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1273), .B1(new_n1277), .B2(new_n1261), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(G2897), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1269), .A2(new_n1239), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n830), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1269), .A2(new_n1239), .A3(G384), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1279), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1275), .B(new_n1276), .C1(new_n1278), .C2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1264), .B1(new_n1278), .B2(new_n1272), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1258), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1254), .A2(new_n1257), .A3(new_n1276), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1263), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1274), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT63), .B1(new_n1278), .B2(new_n1286), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1278), .A2(new_n1272), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1296), .ZN(G405));
  AND3_X1   g1097(.A1(new_n1254), .A2(new_n1257), .A3(new_n1272), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1272), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(G375), .B(new_n1262), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1300), .B(new_n1301), .ZN(G402));
endmodule


