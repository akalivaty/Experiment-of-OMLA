//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n220), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT93), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n224), .A3(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT95), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n216), .B2(new_n217), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT95), .A2(G29gat), .A3(G36gat), .ZN(new_n230));
  AND4_X1   g029(.A1(new_n220), .A2(new_n229), .A3(new_n218), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n214), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT94), .B1(new_n213), .B2(new_n214), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT94), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n210), .A2(new_n212), .A3(new_n234), .A4(KEYINPUT15), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n226), .A2(new_n227), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n227), .B1(new_n226), .B2(new_n236), .ZN(new_n239));
  OAI211_X1 g038(.A(KEYINPUT96), .B(new_n208), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n206), .A2(new_n207), .ZN(new_n241));
  INV_X1    g040(.A(new_n239), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(new_n208), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n240), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(KEYINPUT18), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT97), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n241), .B(new_n245), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n249), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n248), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n249), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n249), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n208), .B1(new_n238), .B2(new_n239), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT96), .B1(new_n241), .B2(new_n245), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n240), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT18), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G141gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G197gat), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT11), .B(G169gat), .Z(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(KEYINPUT12), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n255), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT97), .B1(new_n262), .B2(KEYINPUT18), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n252), .A2(KEYINPUT98), .A3(new_n255), .A4(new_n256), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n263), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n268), .B(KEYINPUT92), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT26), .ZN(new_n284));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n283), .B2(new_n284), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n290), .A2(KEYINPUT28), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT28), .B1(new_n290), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n285), .B1(new_n287), .B2(KEYINPUT24), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n297), .A2(new_n281), .A3(new_n282), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT24), .A3(new_n287), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n295), .B1(new_n299), .B2(new_n298), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT25), .B1(new_n306), .B2(new_n302), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n294), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n309), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G197gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G204gat), .ZN(new_n315));
  INV_X1    g114(.A(G204gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G197gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT22), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G211gat), .ZN(new_n324));
  INV_X1    g123(.A(G218gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n320), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n319), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(KEYINPUT72), .A3(new_n320), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n323), .A2(new_n329), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n315), .B(new_n317), .C1(new_n330), .C2(new_n319), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n330), .A2(new_n319), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n328), .B(new_n327), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n311), .A2(new_n313), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n310), .A2(KEYINPUT74), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n308), .A2(new_n341), .A3(new_n309), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n303), .A2(new_n304), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n302), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n347), .B2(new_n294), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n348), .B2(new_n309), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n337), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n339), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT75), .ZN(new_n355));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  AOI21_X1  g156(.A(new_n280), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n343), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n350), .A2(new_n349), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n280), .B(new_n357), .C1(new_n361), .C2(new_n338), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n360), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n338), .B1(new_n365), .B2(new_n337), .ZN(new_n366));
  INV_X1    g165(.A(new_n357), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR4_X1   g167(.A1(new_n361), .A2(new_n338), .A3(KEYINPUT30), .A4(new_n357), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n358), .A2(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT35), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT64), .ZN(new_n373));
  INV_X1    g172(.A(G127gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(G134gat), .ZN(new_n375));
  INV_X1    g174(.A(G134gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G127gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(G127gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(G134gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT65), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  NAND2_X1  g185(.A1(G113gat), .A2(G120gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT64), .ZN(new_n390));
  AND2_X1   g189(.A1(G113gat), .A2(G120gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(G113gat), .A2(G120gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n381), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G141gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G148gat), .ZN(new_n397));
  INV_X1    g196(.A(G148gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G141gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n397), .A2(new_n399), .B1(KEYINPUT2), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NOR2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT77), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G155gat), .ZN(new_n405));
  INV_X1    g204(.A(G162gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n400), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n401), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n400), .ZN(new_n411));
  XNOR2_X1  g210(.A(G141gat), .B(G148gat), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n400), .A2(KEYINPUT2), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT77), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n391), .A2(new_n392), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n386), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT1), .B1(new_n420), .B2(new_n381), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n378), .C1(new_n421), .C2(new_n390), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n414), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT66), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n389), .B2(new_n394), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT64), .B1(new_n379), .B2(new_n380), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT1), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n417), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT64), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT65), .B1(new_n385), .B2(new_n387), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(KEYINPUT1), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT66), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n433), .A2(new_n440), .A3(KEYINPUT4), .A4(new_n423), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n422), .B1(new_n415), .B2(KEYINPUT3), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT3), .B1(new_n410), .B2(new_n414), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n427), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n431), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n441), .A2(new_n443), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n410), .A2(new_n414), .A3(KEYINPUT3), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n395), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n426), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT78), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n430), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n422), .A2(KEYINPUT4), .A3(new_n423), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n433), .A2(new_n423), .A3(new_n440), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n459), .B2(KEYINPUT4), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G1gat), .B(G29gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G57gat), .B(G85gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n462), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n448), .A2(new_n431), .A3(new_n441), .A4(new_n443), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT78), .B1(new_n450), .B2(new_n453), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n429), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n460), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT6), .B(new_n468), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT81), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n467), .A3(new_n461), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n371), .A2(new_n372), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(KEYINPUT83), .A2(G228gat), .A3(G233gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n337), .B1(new_n446), .B2(KEYINPUT29), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n333), .A2(new_n312), .A3(new_n336), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n423), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n486), .B(new_n487), .C1(new_n489), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n415), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n485), .A3(new_n484), .A4(new_n488), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G22gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G78gat), .B(G106gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(new_n209), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n501), .B(new_n502), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n493), .A2(new_n496), .A3(G22gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(G22gat), .B1(new_n493), .B2(new_n496), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT84), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n507), .B1(new_n512), .B2(new_n503), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n505), .B1(new_n510), .B2(KEYINPUT84), .ZN(new_n514));
  AOI211_X1 g313(.A(new_n508), .B(G22gat), .C1(new_n493), .C2(new_n496), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n507), .B(new_n503), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n506), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n308), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n433), .A2(new_n440), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n294), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G227gat), .ZN(new_n526));
  INV_X1    g325(.A(G233gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n522), .A2(KEYINPUT67), .A3(new_n347), .A4(new_n294), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G43gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT68), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(KEYINPUT68), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT33), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(KEYINPUT32), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n530), .A2(new_n539), .A3(KEYINPUT32), .A4(new_n536), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n530), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n533), .B1(new_n530), .B2(KEYINPUT32), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n538), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n525), .A2(new_n529), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n526), .B2(new_n527), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n544), .A2(new_n548), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n519), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n538), .A2(new_n540), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n542), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n546), .B(KEYINPUT34), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n549), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n483), .A2(new_n518), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n481), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT80), .A4(new_n480), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n370), .B1(new_n565), .B2(new_n477), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT85), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n516), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n570), .A3(new_n548), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n556), .B1(new_n544), .B2(KEYINPUT70), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n569), .A2(new_n506), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g372(.A(new_n561), .B(new_n372), .C1(new_n566), .C2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT6), .B1(new_n462), .B2(new_n468), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT80), .B1(new_n575), .B2(new_n478), .ZN(new_n576));
  INV_X1    g375(.A(new_n564), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n477), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n571), .A2(new_n572), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n371), .A3(new_n579), .A4(new_n518), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT91), .B1(new_n580), .B2(KEYINPUT35), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n560), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT36), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n557), .A2(new_n584), .A3(new_n549), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT86), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n587), .B(new_n588), .C1(new_n566), .C2(new_n518), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n518), .B1(new_n578), .B2(new_n371), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT86), .B1(new_n590), .B2(new_n586), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT39), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n425), .A2(new_n427), .ZN(new_n593));
  OAI221_X1 g392(.A(new_n457), .B1(new_n446), .B2(new_n452), .C1(new_n459), .C2(KEYINPUT4), .ZN(new_n594));
  AOI211_X1 g393(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n427), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT87), .B(KEYINPUT39), .Z(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n427), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n467), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n595), .B2(new_n598), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n370), .A2(new_n479), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n353), .A2(KEYINPUT37), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n604));
  OAI21_X1  g403(.A(new_n357), .B1(new_n353), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT38), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(KEYINPUT38), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n365), .A2(new_n337), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT88), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT88), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n311), .A2(new_n313), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n352), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n609), .B(KEYINPUT37), .C1(new_n608), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n606), .B(new_n614), .C1(new_n353), .C2(new_n357), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n602), .B(new_n518), .C1(new_n615), .C2(new_n482), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n589), .A2(new_n591), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n279), .B1(new_n582), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G57gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(G64gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(G64gat), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(KEYINPUT100), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(KEYINPUT100), .B2(new_n622), .ZN(new_n624));
  NOR2_X1   g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT9), .ZN(new_n626));
  NAND2_X1  g425(.A1(G71gat), .A2(G78gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n622), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n630), .A2(new_n621), .B1(new_n631), .B2(KEYINPUT9), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n625), .B1(new_n631), .B2(new_n627), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n632), .B(new_n633), .C1(new_n631), .C2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(KEYINPUT21), .ZN(new_n637));
  AND2_X1   g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G127gat), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n241), .B1(KEYINPUT21), .B2(new_n636), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n405), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n641), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n640), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(G85gat), .A3(G92gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT7), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT102), .B(G85gat), .Z(new_n656));
  XOR2_X1   g455(.A(KEYINPUT103), .B(G92gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G99gat), .A2(G106gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT8), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G99gat), .B(G106gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n661), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT104), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n661), .B(new_n662), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n665), .B(new_n668), .C1(new_n239), .C2(new_n238), .ZN(new_n669));
  AND2_X1   g468(.A1(G232gat), .A2(G233gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n666), .A2(new_n245), .B1(KEYINPUT41), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT105), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n669), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(G134gat), .B(G162gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n670), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G190gat), .B(G218gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n677), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n673), .A2(new_n675), .A3(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n678), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n681), .B1(new_n678), .B2(new_n683), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(G230gat), .A2(G233gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n664), .A2(new_n635), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n636), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n666), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n689), .A2(new_n690), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  XNOR2_X1  g495(.A(G120gat), .B(G148gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(G176gat), .B(G204gat), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n697), .B(new_n698), .Z(new_n699));
  OR2_X1    g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n694), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(new_n688), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n652), .A2(new_n686), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n619), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n578), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(G1gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1324gat));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n370), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT16), .B(G8gat), .Z(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT107), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(G8gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(KEYINPUT42), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(new_n707), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n720), .B2(new_n587), .ZN(new_n721));
  INV_X1    g520(.A(new_n559), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(G15gat), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n720), .B2(new_n723), .ZN(G1326gat));
  INV_X1    g523(.A(new_n518), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  INV_X1    g527(.A(new_n652), .ZN(new_n729));
  INV_X1    g528(.A(new_n686), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(new_n705), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n279), .B(new_n731), .C1(new_n582), .C2(new_n617), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n216), .A3(new_n708), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT45), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n686), .A2(KEYINPUT44), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n582), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n590), .A2(new_n586), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n616), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n582), .B2(new_n736), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n735), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n582), .A2(new_n617), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n730), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n705), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n279), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n746), .A2(new_n708), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n734), .B1(new_n749), .B2(new_n216), .ZN(G1328gat));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n371), .A2(G36gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n732), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n731), .ZN(new_n754));
  AND4_X1   g553(.A1(new_n751), .A2(new_n618), .A3(new_n754), .A4(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT46), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT110), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n753), .A2(new_n755), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n735), .ZN(new_n761));
  INV_X1    g560(.A(new_n740), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n580), .A2(KEYINPUT35), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n561), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n580), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n722), .A2(new_n725), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n483), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n767), .B2(KEYINPUT108), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n761), .B1(new_n768), .B2(new_n737), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n743), .B2(new_n730), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n370), .B(new_n748), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G36gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(KEYINPUT46), .C1(new_n753), .C2(new_n755), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n757), .A2(new_n760), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT111), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n759), .A2(new_n758), .B1(new_n772), .B2(G36gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n778), .A2(new_n779), .A3(new_n757), .A4(new_n775), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1329gat));
  NAND3_X1  g580(.A1(new_n732), .A2(new_n211), .A3(new_n559), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n746), .A2(new_n586), .A3(new_n748), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(G43gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n785), .B(new_n788), .ZN(G1330gat));
  NAND3_X1  g588(.A1(new_n746), .A2(new_n725), .A3(new_n748), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G50gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n732), .A2(new_n209), .A3(new_n725), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n791), .B(new_n792), .C1(new_n794), .C2(KEYINPUT48), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1331gat));
  NAND2_X1  g598(.A1(new_n279), .A2(new_n704), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n800), .A2(new_n729), .A3(new_n730), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n738), .B2(new_n741), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(new_n578), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G57gat), .ZN(G1332gat));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(KEYINPUT114), .B(new_n801), .C1(new_n738), .C2(new_n741), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n370), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT49), .B(G64gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n806), .A2(new_n370), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n810), .B1(new_n809), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1333gat));
  NAND4_X1  g614(.A1(new_n806), .A2(G71gat), .A3(new_n586), .A4(new_n807), .ZN(new_n816));
  INV_X1    g615(.A(G71gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n802), .B2(new_n722), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g619(.A1(new_n806), .A2(new_n725), .A3(new_n807), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g621(.A1(new_n800), .A2(new_n652), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n746), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n708), .ZN(new_n825));
  INV_X1    g624(.A(new_n279), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n652), .A3(new_n686), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n768), .B2(new_n737), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT51), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n829), .A2(KEYINPUT51), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(KEYINPUT116), .A3(KEYINPUT51), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n708), .A2(new_n656), .A3(new_n704), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT117), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n825), .A2(new_n656), .B1(new_n835), .B2(new_n837), .ZN(G1336gat));
  NAND3_X1  g637(.A1(new_n746), .A2(new_n370), .A3(new_n823), .ZN(new_n839));
  INV_X1    g638(.A(new_n657), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n371), .A2(new_n705), .A3(G92gat), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n835), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n839), .A2(new_n840), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n833), .B2(new_n830), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT52), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(G1337gat));
  NAND2_X1  g647(.A1(new_n824), .A2(new_n586), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT118), .B(G99gat), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n722), .A2(new_n705), .A3(new_n850), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n835), .B2(new_n852), .ZN(G1338gat));
  NAND3_X1  g652(.A1(new_n746), .A2(new_n725), .A3(new_n823), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT53), .B1(new_n854), .B2(G106gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n518), .A2(new_n705), .A3(G106gat), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n855), .B1(new_n835), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n854), .A2(G106gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n833), .B2(new_n830), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT53), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(G1339gat));
  OR2_X1    g661(.A1(new_n706), .A2(new_n826), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n692), .A2(new_n693), .A3(new_n688), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n701), .A2(KEYINPUT54), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n699), .B1(new_n694), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(KEYINPUT55), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(new_n703), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n867), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n869), .B(new_n872), .C1(new_n684), .C2(new_n685), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n257), .A2(new_n270), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n248), .A2(new_n249), .B1(new_n253), .B2(new_n254), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n267), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n704), .A3(new_n876), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n869), .A2(new_n872), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n279), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n881), .B2(new_n686), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n863), .B1(new_n882), .B2(new_n652), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n766), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n578), .A2(new_n370), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n279), .A2(new_n383), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n883), .A2(new_n708), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(new_n573), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n371), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n383), .B1(new_n893), .B2(new_n279), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT120), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n890), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1340gat));
  NAND3_X1  g698(.A1(new_n888), .A2(G120gat), .A3(new_n704), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n384), .B1(new_n893), .B2(new_n705), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(G1341gat));
  XNOR2_X1  g701(.A(new_n886), .B(KEYINPUT119), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n374), .A3(new_n729), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n729), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(G127gat), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT121), .B1(new_n893), .B2(new_n729), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(G1342gat));
  NOR2_X1   g707(.A1(new_n686), .A2(new_n370), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n376), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT56), .Z(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n903), .B2(new_n686), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1343gat));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n883), .B2(new_n725), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n883), .A2(KEYINPUT57), .A3(new_n725), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n586), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n885), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n918), .B2(new_n279), .ZN(new_n919));
  AND4_X1   g718(.A1(new_n708), .A2(new_n883), .A3(new_n725), .A4(new_n587), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n920), .A2(new_n371), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n396), .A3(new_n826), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(KEYINPUT58), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1344gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n398), .A3(new_n704), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n705), .B1(new_n915), .B2(new_n916), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n586), .A2(new_n578), .A3(new_n370), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n398), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n930), .B(KEYINPUT122), .Z(new_n932));
  AND2_X1   g731(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n934));
  OAI221_X1 g733(.A(new_n928), .B1(new_n931), .B2(KEYINPUT59), .C1(new_n933), .C2(new_n934), .ZN(G1345gat));
  OAI21_X1  g734(.A(G155gat), .B1(new_n918), .B2(new_n729), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n405), .A3(new_n652), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT123), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(G162gat), .B1(new_n918), .B2(new_n686), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n920), .A2(new_n406), .A3(new_n909), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n708), .A2(new_n371), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n884), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n884), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(new_n281), .A3(new_n279), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n883), .A2(new_n578), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(new_n370), .A3(new_n573), .ZN(new_n954));
  AOI21_X1  g753(.A(G169gat), .B1(new_n954), .B2(new_n826), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n952), .A2(new_n955), .ZN(G1348gat));
  OAI21_X1  g755(.A(G176gat), .B1(new_n951), .B2(new_n705), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n954), .A2(new_n282), .A3(new_n704), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n951), .B2(new_n729), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(new_n290), .A3(new_n652), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n954), .A2(new_n291), .A3(new_n730), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n730), .A3(new_n950), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n968), .A2(new_n969), .A3(G190gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n968), .B2(G190gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  NOR3_X1   g771(.A1(new_n586), .A2(new_n371), .A3(new_n518), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n953), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(G197gat), .A3(new_n279), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT125), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n883), .A2(KEYINPUT57), .A3(new_n725), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n587), .B(new_n946), .C1(new_n977), .C2(new_n914), .ZN(new_n978));
  OAI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n279), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(G1352gat));
  INV_X1    g779(.A(KEYINPUT62), .ZN(new_n981));
  INV_X1    g780(.A(new_n974), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n982), .A2(new_n316), .A3(new_n704), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n981), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n986), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n988), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n989));
  OAI21_X1  g788(.A(G204gat), .B1(new_n978), .B2(new_n705), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n982), .A2(new_n324), .A3(new_n652), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n978), .A2(new_n729), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n324), .B1(new_n993), .B2(KEYINPUT127), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n978), .B2(new_n729), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n917), .A2(KEYINPUT127), .A3(new_n652), .A4(new_n946), .ZN(new_n998));
  AND4_X1   g797(.A1(KEYINPUT63), .A2(new_n998), .A3(G211gat), .A4(new_n996), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(G1354gat));
  OAI21_X1  g799(.A(G218gat), .B1(new_n978), .B2(new_n686), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n982), .A2(new_n325), .A3(new_n730), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1355gat));
endmodule


