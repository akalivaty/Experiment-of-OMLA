//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n567, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT69), .B(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n462), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(KEYINPUT69), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n479), .A2(new_n482), .A3(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(G124), .B2(new_n496), .ZN(G162));
  NAND2_X1  g072(.A1(new_n470), .A2(G102), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n492), .A2(new_n480), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G114), .A2(G2104), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n480), .B2(G126), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n498), .B(new_n502), .C1(new_n505), .C2(new_n483), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT4), .B1(new_n468), .B2(G138), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .A3(G62), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n511), .B(new_n513), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n528), .A3(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(G543), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n522), .A2(new_n534), .ZN(G166));
  AND2_X1   g110(.A1(new_n527), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  INV_X1    g112(.A(new_n524), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT6), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n510), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n537), .A2(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n536), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n514), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(G52), .B2(new_n540), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n514), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(G43), .B2(new_n540), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT74), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT75), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G188));
  XNOR2_X1  g143(.A(new_n518), .B(KEYINPUT77), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G65), .ZN(new_n570));
  INV_X1    g145(.A(G78), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n510), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(G91), .B2(new_n536), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n533), .A2(KEYINPUT76), .A3(new_n574), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT9), .Z(new_n576));
  NAND2_X1  g151(.A1(new_n573), .A2(new_n576), .ZN(G299));
  OAI221_X1 g152(.A(new_n521), .B1(new_n532), .B2(new_n533), .C1(new_n531), .C2(new_n530), .ZN(G303));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n514), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n540), .B2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n527), .A2(G87), .A3(new_n529), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n511), .A2(new_n513), .A3(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n540), .B2(G48), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n527), .A2(G86), .A3(new_n529), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n540), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n591), .B2(new_n592), .C1(new_n530), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n533), .A2(KEYINPUT78), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n533), .A2(KEYINPUT78), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n596), .A2(G54), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n530), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n536), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n569), .A2(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n605), .B2(new_n510), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n605), .A2(new_n510), .A3(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n595), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n595), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  XNOR2_X1  g191(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n480), .A2(new_n470), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  OAI221_X1 g202(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n492), .C2(G111), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n628), .B1(new_n495), .B2(new_n629), .C1(new_n630), .C2(new_n484), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT83), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2443), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT17), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n652), .A2(new_n657), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  XOR2_X1   g237(.A(new_n652), .B(KEYINPUT85), .Z(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n662), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n669), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  AOI22_X1  g250(.A1(new_n673), .A2(KEYINPUT20), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n669), .A3(new_n672), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n676), .B(new_n678), .C1(KEYINPUT20), .C2(new_n673), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT86), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G26), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n496), .A2(G128), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n485), .A2(G140), .ZN(new_n690));
  OAI221_X1 g265(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n492), .C2(G116), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n688), .B1(new_n693), .B2(new_n687), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n688), .B(new_n694), .S(KEYINPUT28), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT93), .B(G2067), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n492), .A2(G103), .A3(G2104), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT25), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n485), .A2(G139), .ZN(new_n700));
  AOI22_X1  g275(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n700), .C1(new_n492), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G33), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G2072), .Z(new_n704));
  NAND2_X1  g279(.A1(G171), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G5), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1961), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT95), .Z(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT94), .B1(new_n470), .B2(G105), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n470), .A2(KEYINPUT94), .A3(G105), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n496), .A2(G129), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G141), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G29), .B2(G32), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G168), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G16), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  NAND2_X1  g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n729), .A2(new_n730), .A3(G29), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n726), .A2(new_n727), .B1(G2084), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n704), .A2(new_n708), .A3(new_n724), .A4(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n697), .B(new_n736), .C1(new_n737), .C2(new_n733), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n726), .A2(new_n727), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT97), .Z(new_n740));
  NOR2_X1   g315(.A1(new_n706), .A2(new_n707), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT99), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n687), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n687), .ZN(new_n744));
  MUX2_X1   g319(.A(new_n743), .B(new_n744), .S(KEYINPUT100), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2078), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  INV_X1    g322(.A(G28), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n749), .A2(new_n750), .A3(new_n687), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n747), .B(new_n751), .C1(new_n631), .C2(new_n687), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n740), .A2(new_n742), .A3(new_n746), .A4(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n721), .A2(new_n723), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n611), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT91), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1348), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n738), .A2(new_n754), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G16), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n761), .A2(KEYINPUT92), .A3(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n561), .B2(new_n761), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT92), .B1(new_n761), .B2(G19), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  OAI21_X1  g341(.A(KEYINPUT23), .B1(new_n615), .B2(new_n761), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n761), .A2(G20), .ZN(new_n768));
  MUX2_X1   g343(.A(KEYINPUT23), .B(new_n767), .S(new_n768), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n760), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G23), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n581), .A2(new_n582), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(G288), .A2(KEYINPUT88), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G16), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XOR2_X1   g354(.A(new_n778), .B(new_n779), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n761), .A2(G22), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G166), .B2(new_n761), .ZN(new_n782));
  INV_X1    g357(.A(G1971), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n761), .A2(G6), .ZN(new_n785));
  INV_X1    g360(.A(G305), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n761), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT32), .B(G1981), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n780), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT89), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n687), .A2(G25), .ZN(new_n793));
  INV_X1    g368(.A(G119), .ZN(new_n794));
  OR3_X1    g369(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT87), .B1(new_n495), .B2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n795), .A2(new_n796), .B1(G131), .B2(new_n485), .ZN(new_n797));
  OAI221_X1 g372(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n492), .C2(G107), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n793), .B1(new_n800), .B2(new_n687), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT35), .B(G1991), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n806));
  OR2_X1    g381(.A1(G16), .A2(G24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G290), .B2(new_n761), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n792), .A2(new_n804), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT36), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n687), .A2(G35), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G162), .B2(new_n687), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT29), .B(G2090), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n792), .A2(KEYINPUT36), .A3(new_n804), .A4(new_n812), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n771), .A2(new_n815), .A3(new_n819), .A4(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  NAND2_X1  g397(.A1(new_n536), .A2(G93), .ZN(new_n823));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n514), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n826), .A2(G651), .B1(G55), .B2(new_n540), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT102), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n611), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n561), .A2(new_n828), .ZN(new_n834));
  INV_X1    g409(.A(new_n828), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(new_n560), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n833), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n839), .B2(KEYINPUT101), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(KEYINPUT101), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n831), .B1(new_n841), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n631), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n799), .B(new_n718), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n625), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI221_X1 g427(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n492), .C2(G118), .ZN(new_n853));
  INV_X1    g428(.A(G142), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n484), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G130), .B2(new_n496), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n702), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n692), .B(G164), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n857), .B(new_n858), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n850), .A2(new_n861), .A3(new_n851), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n777), .B(G290), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G166), .B(KEYINPUT105), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n786), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n868), .A3(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n837), .B(new_n620), .Z(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n610), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n573), .A2(new_n603), .A3(new_n576), .A4(new_n609), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n837), .B(new_n620), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n882));
  AND2_X1   g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n880), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n874), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  INV_X1    g466(.A(new_n874), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G868), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n835), .A2(G868), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n866), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g473(.A(KEYINPUT107), .B(new_n896), .C1(new_n894), .C2(G868), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G295));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n897), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n874), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n883), .A2(new_n884), .ZN(new_n904));
  XNOR2_X1  g479(.A(G286), .B(G301), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n837), .B(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n879), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n874), .B(new_n902), .C1(new_n909), .C2(new_n907), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n863), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n878), .A2(new_n916), .A3(KEYINPUT41), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n878), .B2(KEYINPUT41), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n878), .A2(new_n882), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(KEYINPUT110), .B(new_n908), .C1(new_n920), .C2(new_n906), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(new_n874), .C1(KEYINPUT110), .C2(new_n908), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n892), .A2(new_n910), .ZN(new_n923));
  AND4_X1   g498(.A1(KEYINPUT43), .A2(new_n922), .A3(new_n863), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT44), .B1(new_n915), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n914), .A4(new_n863), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n506), .B2(new_n507), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n476), .A2(new_n469), .A3(G40), .A4(new_n471), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n718), .B(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n692), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n802), .B2(new_n799), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n800), .A2(new_n803), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G290), .B(new_n809), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(G8), .B1(new_n933), .B2(new_n936), .ZN(new_n949));
  NAND2_X1  g524(.A1(G305), .A2(G1981), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n587), .A2(new_n588), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT113), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT49), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n950), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n949), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1976), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n773), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n949), .B1(new_n966), .B2(new_n953), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n936), .B1(new_n933), .B2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n932), .C1(new_n506), .C2(new_n507), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT111), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n492), .A2(new_n480), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n499), .B1(new_n972), .B2(new_n500), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n503), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G2105), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n976), .A3(new_n498), .A4(new_n502), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n969), .A4(new_n932), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT118), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n968), .A2(new_n971), .A3(new_n982), .A4(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n707), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n985));
  INV_X1    g560(.A(new_n936), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n977), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n935), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n988), .B2(G2078), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n935), .A2(new_n987), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(KEYINPUT53), .A3(new_n991), .A4(new_n986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G171), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(G168), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n988), .A2(new_n727), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n968), .A2(new_n971), .A3(new_n737), .A4(new_n979), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(G8), .ZN(new_n1004));
  INV_X1    g579(.A(new_n997), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1007), .A2(new_n997), .A3(new_n999), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1009), .A3(new_n997), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n1003), .B2(new_n997), .ZN(new_n1012));
  OAI22_X1  g587(.A1(new_n1006), .A2(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n994), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n777), .A2(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n965), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n963), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n965), .B1(new_n775), .B2(new_n776), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT52), .B1(new_n1018), .B2(new_n949), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n964), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1021));
  NAND3_X1  g596(.A1(G303), .A2(G8), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n522), .B2(new_n534), .ZN(new_n1023));
  NAND2_X1  g598(.A1(KEYINPUT112), .A2(KEYINPUT55), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n933), .A2(KEYINPUT50), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1028), .A2(new_n986), .A3(new_n970), .ZN(new_n1029));
  INV_X1    g604(.A(G2090), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1029), .A2(new_n1030), .B1(new_n988), .B2(new_n783), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1031), .B2(new_n996), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n988), .A2(new_n783), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n968), .A2(new_n971), .A3(new_n1030), .A4(new_n979), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n996), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1026), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1020), .A2(new_n1032), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1004), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n999), .B1(new_n1007), .B2(new_n997), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1003), .A2(new_n997), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT121), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1038), .A2(new_n1039), .B1(new_n1041), .B2(new_n1010), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n967), .B1(new_n1014), .B2(new_n1044), .ZN(new_n1045));
  AOI221_X4 g620(.A(new_n996), .B1(new_n1022), .B2(new_n1025), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1020), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n996), .B(G286), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1020), .A2(new_n1036), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT63), .B1(new_n1035), .B2(new_n1026), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n964), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1046), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1057), .B2(new_n1027), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1054), .A2(KEYINPUT115), .A3(new_n1058), .A4(new_n1049), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1020), .A2(new_n1032), .A3(new_n1036), .A4(new_n1049), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT114), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n1055), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1045), .A2(new_n1047), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1348), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n981), .A2(new_n1068), .A3(new_n983), .ZN(new_n1069));
  INV_X1    g644(.A(new_n933), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n941), .A3(new_n986), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT117), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n611), .A2(KEYINPUT120), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n610), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(new_n610), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n935), .A2(new_n986), .A3(new_n987), .A4(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n968), .A2(new_n970), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G299), .B(KEYINPUT57), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1083), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1086), .A2(KEYINPUT119), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n933), .B2(new_n936), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n988), .B2(G1996), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n561), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT59), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1082), .A2(new_n1095), .A3(new_n1101), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1100), .A2(new_n611), .A3(new_n1078), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1108), .A2(new_n1099), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n475), .B(KEYINPUT123), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n985), .B(new_n472), .C1(new_n1111), .C2(new_n467), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n990), .A2(G40), .A3(new_n991), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n984), .A2(new_n989), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n984), .A2(KEYINPUT124), .A3(new_n989), .A4(new_n1113), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(G171), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n984), .A2(G301), .A3(new_n989), .A4(new_n992), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(KEYINPUT54), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT125), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1118), .A2(new_n1123), .A3(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n994), .B1(G171), .B2(new_n1114), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1037), .B(new_n1042), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1110), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n948), .B1(new_n1067), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n937), .A2(new_n939), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT46), .Z(new_n1132));
  AOI21_X1  g707(.A(new_n938), .B1(new_n942), .B2(new_n719), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT47), .Z(new_n1135));
  NOR3_X1   g710(.A1(new_n938), .A2(G1986), .A3(G290), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT48), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n946), .B2(new_n938), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n945), .B(KEYINPUT126), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1139), .A2(new_n943), .B1(G2067), .B2(new_n692), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n937), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT127), .B1(new_n1130), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1142), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1014), .A2(new_n1044), .ZN(new_n1146));
  INV_X1    g721(.A(new_n967), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1066), .A2(new_n1146), .A3(new_n1047), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1127), .A2(new_n1126), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1037), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1013), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1151), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1110), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1144), .B(new_n1145), .C1(new_n1153), .C2(new_n948), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1143), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g730(.A1(new_n864), .A2(new_n649), .A3(new_n666), .ZN(new_n1157));
  INV_X1    g731(.A(G319), .ZN(new_n1158));
  NOR2_X1   g732(.A1(G229), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n928), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


