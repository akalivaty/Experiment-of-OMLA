//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n809, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT14), .B(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(KEYINPUT96), .A3(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT96), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  INV_X1    g017(.A(new_n207), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n203), .B2(new_n204), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n212), .B1(new_n221), .B2(new_n211), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n202), .B1(new_n222), .B2(KEYINPUT97), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n220), .A2(new_n210), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n209), .A2(new_n217), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n208), .B1(new_n225), .B2(new_n216), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n226), .B2(new_n210), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT97), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(KEYINPUT98), .C1(G1gat), .C2(new_n231), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n237), .A2(KEYINPUT99), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(KEYINPUT99), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n237), .A2(new_n222), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .A4(new_n242), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n237), .B(new_n222), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n241), .B(KEYINPUT13), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT95), .ZN(new_n251));
  XNOR2_X1  g050(.A(G169gat), .B(G197gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT94), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G113gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n255));
  INV_X1    g054(.A(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n254), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n250), .A2(KEYINPUT95), .A3(new_n259), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n265), .A2(G169gat), .A3(G176gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n264), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT23), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT65), .A3(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT25), .B1(new_n275), .B2(KEYINPUT23), .ZN(new_n276));
  OR2_X1    g075(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n276), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n265), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n272), .A2(new_n296), .A3(new_n267), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n288), .A2(new_n290), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G226gat), .ZN(new_n301));
  INV_X1    g100(.A(G233gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n305), .A2(new_n281), .ZN(new_n306));
  INV_X1    g105(.A(new_n275), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n267), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G183gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n315), .A2(new_n277), .A3(new_n279), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n278), .A2(KEYINPUT27), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n314), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n277), .A2(new_n279), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT28), .A3(new_n313), .A4(new_n317), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n310), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n300), .A2(new_n304), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n330), .B(new_n331), .Z(new_n332));
  AOI21_X1  g131(.A(new_n298), .B1(new_n287), .B2(KEYINPUT67), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n322), .B1(new_n333), .B2(new_n290), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n303), .A2(KEYINPUT29), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n324), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n300), .A2(new_n323), .ZN(new_n338));
  INV_X1    g137(.A(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n332), .A4(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n332), .B(KEYINPUT75), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n340), .B2(new_n324), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n345), .B1(new_n337), .B2(new_n342), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT30), .A3(new_n349), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n343), .A2(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n359));
  INV_X1    g158(.A(new_n349), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G148gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n256), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT78), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT2), .ZN(new_n373));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n369), .A2(new_n371), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G155gat), .ZN(new_n377));
  INV_X1    g176(.A(G155gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT80), .B(G162gat), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n370), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n369), .A2(new_n377), .A3(new_n379), .A4(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389));
  INV_X1    g188(.A(G113gat), .ZN(new_n390));
  INV_X1    g189(.A(G120gat), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT1), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(KEYINPUT69), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G113gat), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n391), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(G113gat), .B2(G120gat), .ZN(new_n399));
  AND2_X1   g198(.A1(G113gat), .A2(G120gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n393), .A2(new_n397), .B1(new_n401), .B2(new_n389), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n388), .A2(new_n402), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n377), .A2(new_n369), .A3(new_n379), .A4(new_n374), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n376), .ZN(new_n406));
  NAND2_X1  g205(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n382), .A2(new_n383), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n408), .B2(new_n370), .ZN(new_n409));
  INV_X1    g208(.A(G134gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G127gat), .ZN(new_n411));
  INV_X1    g210(.A(G127gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G134gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n399), .B2(new_n400), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT69), .B(G113gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n392), .B(new_n389), .C1(new_n416), .C2(new_n391), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n409), .A2(new_n381), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n367), .B1(new_n403), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n422));
  AND2_X1   g221(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n423));
  AND2_X1   g222(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(KEYINPUT80), .A2(G162gat), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n422), .A2(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT2), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n427), .A2(new_n404), .B1(new_n380), .B2(new_n375), .ZN(new_n428));
  INV_X1    g227(.A(new_n397), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n399), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n392), .B1(new_n390), .B2(new_n391), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n429), .A2(new_n430), .B1(new_n431), .B2(new_n414), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n388), .A2(new_n402), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(KEYINPUT81), .A3(new_n367), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n432), .B1(new_n428), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n367), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n417), .A2(KEYINPUT70), .A3(new_n415), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT70), .B1(new_n417), .B2(new_n415), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n428), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(KEYINPUT5), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n402), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n417), .A2(KEYINPUT70), .A3(new_n415), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n428), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n442), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n409), .A2(new_n438), .A3(new_n381), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n402), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n366), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n365), .B1(new_n449), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n456), .A2(new_n460), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n453), .A2(KEYINPUT4), .ZN(new_n467));
  INV_X1    g266(.A(new_n447), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n469), .B2(new_n441), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n466), .B1(new_n470), .B2(new_n437), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n471), .B2(new_n365), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n463), .B1(new_n472), .B2(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n365), .A3(new_n461), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n464), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n421), .A2(new_n436), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n447), .B1(KEYINPUT4), .B2(new_n453), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n366), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT5), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n461), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n365), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n465), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n465), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n355), .B(new_n361), .C1(new_n476), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n330), .B(new_n331), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n438), .B1(new_n489), .B2(KEYINPUT29), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n388), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n428), .B2(new_n438), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n332), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G228gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n302), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT86), .B(G22gat), .Z(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n302), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n491), .B(new_n497), .C1(new_n344), .C2(new_n492), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n501));
  XOR2_X1   g300(.A(G78gat), .B(G106gat), .Z(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT31), .B(G50gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n495), .A2(new_n498), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G22gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n504), .B(KEYINPUT85), .ZN(new_n508));
  INV_X1    g307(.A(new_n499), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n496), .B1(new_n495), .B2(new_n498), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  INV_X1    g314(.A(G227gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n302), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n300), .A2(new_n445), .A3(new_n323), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n445), .B1(new_n300), .B2(new_n323), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G15gat), .B(G43gat), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT71), .ZN(new_n522));
  XNOR2_X1  g321(.A(G71gat), .B(G99gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT33), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n527), .A3(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(new_n517), .ZN(new_n529));
  INV_X1    g328(.A(new_n445), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n338), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n334), .A2(new_n445), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n533), .A2(KEYINPUT33), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n529), .A3(new_n532), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT34), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(KEYINPUT34), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n520), .A2(KEYINPUT32), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n520), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n545), .A3(new_n524), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n546), .A2(new_n528), .B1(new_n540), .B2(new_n539), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n515), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n539), .A2(new_n540), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n551), .A2(new_n537), .A3(KEYINPUT73), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n537), .B2(KEYINPUT73), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT36), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g353(.A(KEYINPUT74), .B(new_n515), .C1(new_n542), .C2(new_n547), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n358), .A2(KEYINPUT37), .A3(new_n359), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n345), .A2(KEYINPUT37), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n349), .B1(new_n343), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n343), .A2(new_n559), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n303), .B(new_n322), .C1(new_n333), .C2(new_n290), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n335), .B1(new_n300), .B2(new_n323), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n489), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n344), .B(new_n324), .C1(new_n334), .C2(new_n335), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT89), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n568), .B(new_n489), .C1(new_n563), .C2(new_n564), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(KEYINPUT37), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n349), .A2(KEYINPUT38), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n562), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT90), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n562), .A2(new_n570), .A3(new_n574), .A4(new_n571), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n463), .A2(new_n472), .B1(new_n353), .B2(new_n349), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT91), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT84), .B1(new_n462), .B2(new_n465), .ZN(new_n579));
  NOR4_X1   g378(.A1(new_n471), .A2(new_n484), .A3(new_n365), .A4(new_n464), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n485), .A2(KEYINPUT91), .A3(new_n486), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n561), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n585));
  AOI211_X1 g384(.A(new_n357), .B(new_n345), .C1(new_n337), .C2(new_n342), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n585), .A2(new_n586), .A3(new_n349), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n352), .A2(new_n354), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n458), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n367), .B1(new_n456), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n591), .B(KEYINPUT39), .C1(new_n367), .C2(new_n435), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n367), .C1(new_n456), .C2(new_n590), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT88), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n594), .A2(new_n595), .A3(new_n365), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n594), .B2(new_n365), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n592), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n462), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n599), .B2(new_n598), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n512), .B1(new_n589), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n514), .B(new_n556), .C1(new_n584), .C2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n512), .B1(new_n552), .B2(new_n553), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n488), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n542), .B2(new_n547), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n551), .A2(new_n528), .A3(new_n546), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n537), .A2(new_n541), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(KEYINPUT92), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n463), .A2(new_n472), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n582), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT35), .B1(new_n507), .B2(new_n511), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(new_n589), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n605), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n263), .B1(new_n603), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g427(.A(G99gat), .B(G106gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(G92gat), .ZN(new_n630));
  INV_X1    g429(.A(G85gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n630), .A2(new_n631), .B1(KEYINPUT8), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n628), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n223), .B2(new_n229), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n637), .A2(new_n227), .B1(KEYINPUT41), .B2(new_n618), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n624), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n618), .A2(KEYINPUT41), .ZN(new_n642));
  INV_X1    g441(.A(new_n637), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n222), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n638), .A2(new_n644), .A3(new_n623), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n622), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n624), .A3(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n623), .B1(new_n638), .B2(new_n644), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n621), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT21), .ZN(new_n652));
  INV_X1    g451(.A(G57gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(G64gat), .ZN(new_n654));
  INV_X1    g453(.A(G64gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(G57gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n657), .B2(KEYINPUT100), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G71gat), .B(G78gat), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n656), .A2(KEYINPUT101), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(KEYINPUT101), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n665), .A3(new_n654), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n237), .B(new_n651), .C1(new_n652), .C2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n237), .B1(new_n652), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT103), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n661), .A2(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n673));
  OAI211_X1 g472(.A(G231gat), .B(G233gat), .C1(new_n673), .C2(KEYINPUT21), .ZN(new_n674));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n652), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n676), .A3(new_n412), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n412), .B1(new_n674), .B2(new_n676), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n670), .B(new_n672), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n672), .A2(new_n670), .ZN(new_n681));
  INV_X1    g480(.A(new_n679), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n677), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G155gat), .ZN(new_n686));
  XOR2_X1   g485(.A(G183gat), .B(G211gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n680), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n680), .B2(new_n683), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n650), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n689), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT106), .A3(new_n650), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(G230gat), .A2(G233gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n669), .B1(new_n635), .B2(new_n636), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT10), .ZN(new_n702));
  INV_X1    g501(.A(new_n636), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n673), .A2(new_n703), .A3(new_n634), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n637), .A2(KEYINPUT10), .A3(new_n673), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT107), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n700), .C1(new_n705), .C2(new_n706), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n699), .B1(new_n701), .B2(new_n704), .ZN(new_n712));
  XNOR2_X1  g511(.A(G120gat), .B(G148gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(G176gat), .B(G204gat), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n713), .B(new_n714), .Z(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n707), .B2(new_n712), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n698), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n617), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n476), .A2(new_n487), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G1gat), .ZN(G1324gat));
  INV_X1    g524(.A(new_n589), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n728), .A2(G8gat), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT16), .B(G8gat), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n727), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n728), .B2(new_n729), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n730), .B(new_n733), .C1(new_n734), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g534(.A(new_n722), .ZN(new_n736));
  OAI21_X1  g535(.A(G15gat), .B1(new_n736), .B2(new_n556), .ZN(new_n737));
  INV_X1    g536(.A(new_n611), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(G15gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n736), .B2(new_n739), .ZN(G1326gat));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n513), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT43), .B(G22gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1327gat));
  NOR3_X1   g542(.A1(new_n720), .A2(new_n696), .A3(new_n650), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT109), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n617), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n206), .A3(new_n723), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT45), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750));
  INV_X1    g549(.A(new_n262), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n259), .B1(new_n250), .B2(KEYINPUT95), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n261), .A2(KEYINPUT110), .A3(new_n262), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(new_n696), .A3(new_n720), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n603), .A2(new_n616), .ZN(new_n758));
  INV_X1    g557(.A(new_n650), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n650), .B(new_n762), .C1(new_n603), .C2(new_n616), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n756), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT112), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n766), .B(new_n756), .C1(new_n760), .C2(new_n763), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n765), .A2(new_n723), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n749), .B1(new_n768), .B2(new_n206), .ZN(G1328gat));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n726), .A3(new_n767), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT113), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n765), .A2(new_n772), .A3(new_n726), .A4(new_n767), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(G36gat), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n746), .A2(G36gat), .A3(new_n589), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT46), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1329gat));
  NOR3_X1   g576(.A1(new_n746), .A2(G43gat), .A3(new_n738), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(KEYINPUT114), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n556), .ZN(new_n781));
  NAND2_X1  g580(.A1(KEYINPUT47), .A2(G43gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n556), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n765), .A2(new_n784), .A3(new_n767), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n785), .A2(G43gat), .B1(KEYINPUT114), .B2(new_n778), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g586(.A(G50gat), .B1(new_n764), .B2(new_n512), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n746), .A2(G50gat), .A3(new_n512), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(KEYINPUT48), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n765), .A2(new_n513), .A3(new_n767), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n792), .B2(G50gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n793), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g593(.A(new_n698), .B1(new_n753), .B2(new_n754), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n720), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n603), .B2(new_n616), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n723), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g598(.A(new_n589), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT115), .ZN(new_n802));
  NOR2_X1   g601(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1333gat));
  NAND2_X1  g603(.A1(new_n797), .A2(new_n784), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n738), .A2(G71gat), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n805), .A2(G71gat), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g607(.A1(new_n797), .A2(new_n513), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G78gat), .ZN(G1335gat));
  INV_X1    g609(.A(new_n755), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n696), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n719), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n711), .B2(new_n717), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n760), .B2(new_n763), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT116), .B(new_n816), .C1(new_n760), .C2(new_n763), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n723), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G85gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n758), .A2(new_n759), .A3(new_n812), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n815), .B1(new_n823), .B2(KEYINPUT51), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(KEYINPUT51), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n723), .A2(new_n631), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(G1336gat));
  INV_X1    g626(.A(new_n630), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n817), .B2(new_n589), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n589), .A2(G92gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n829), .B(new_n830), .C1(new_n825), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n825), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n726), .A3(new_n820), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(new_n828), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n833), .B1(new_n836), .B2(new_n830), .ZN(G1337gat));
  INV_X1    g636(.A(G99gat), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n825), .A2(new_n738), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n819), .A2(new_n820), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n556), .A2(new_n838), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(G1338gat));
  OAI21_X1  g641(.A(G106gat), .B1(new_n817), .B2(new_n512), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n512), .A2(G106gat), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n843), .B(new_n844), .C1(new_n825), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n825), .A2(new_n846), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n819), .A2(new_n513), .A3(new_n820), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(G106gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n844), .ZN(G1339gat));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n795), .B2(new_n815), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n694), .A2(new_n697), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n852), .A2(new_n755), .A3(new_n854), .A4(new_n815), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n696), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n705), .A2(new_n706), .A3(new_n700), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n708), .A2(new_n710), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n715), .B1(new_n707), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n858), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n707), .B(KEYINPUT107), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT55), .B(new_n863), .C1(new_n866), .C2(new_n860), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n865), .A2(new_n867), .A3(new_n718), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n753), .A2(new_n754), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n241), .B1(new_n240), .B2(new_n242), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n247), .A2(new_n248), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n258), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n245), .A2(new_n246), .A3(new_n249), .A4(new_n259), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n720), .A2(new_n870), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n873), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n876), .B2(new_n815), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n759), .B1(new_n869), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n865), .A2(new_n867), .A3(new_n718), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n650), .A3(new_n876), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n857), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n513), .B1(new_n856), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n723), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n726), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n738), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n263), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n883), .A2(KEYINPUT119), .A3(new_n887), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G113gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n795), .A2(new_n852), .A3(new_n815), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n755), .A2(new_n854), .A3(new_n815), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT117), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n726), .A2(new_n604), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n723), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n416), .A3(new_n811), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n894), .A2(new_n901), .ZN(G1340gat));
  AOI21_X1  g701(.A(G120gat), .B1(new_n900), .B2(new_n720), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n890), .A2(new_n892), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n815), .A2(new_n391), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(G1341gat));
  AND2_X1   g705(.A1(new_n900), .A2(new_n696), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n908));
  AOI21_X1  g707(.A(G127gat), .B1(new_n907), .B2(KEYINPUT120), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n857), .A2(new_n412), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n908), .A2(new_n909), .B1(new_n904), .B2(new_n910), .ZN(G1342gat));
  NAND3_X1  g710(.A1(new_n900), .A2(new_n410), .A3(new_n759), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(KEYINPUT121), .B2(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g712(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n890), .A2(new_n759), .A3(new_n892), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G134gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n912), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(G1343gat));
  NOR3_X1   g718(.A1(new_n784), .A2(new_n512), .A3(new_n726), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n263), .A2(G141gat), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n898), .A2(new_n723), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n886), .A2(new_n784), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n869), .A2(new_n878), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n650), .ZN(new_n928));
  INV_X1    g727(.A(new_n881), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n696), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n895), .A2(new_n897), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n513), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n720), .A2(KEYINPUT122), .A3(new_n873), .A4(new_n874), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n876), .B2(new_n815), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n935), .B(new_n937), .C1(new_n263), .C2(new_n880), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(new_n650), .ZN(new_n939));
  OAI211_X1 g738(.A(KEYINPUT123), .B(new_n857), .C1(new_n939), .C2(new_n881), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n881), .B1(new_n938), .B2(new_n650), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n696), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n856), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n512), .A2(new_n933), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n263), .B(new_n926), .C1(new_n934), .C2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n924), .B1(new_n947), .B2(new_n256), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT58), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n944), .A2(new_n945), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT57), .B1(new_n898), .B2(new_n513), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n925), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G141gat), .B1(new_n952), .B2(new_n755), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n954), .A2(new_n955), .A3(new_n949), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n948), .A2(new_n949), .B1(new_n953), .B2(new_n956), .ZN(G1344gat));
  AND3_X1   g756(.A1(new_n898), .A2(new_n723), .A3(new_n920), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n368), .A3(new_n720), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n926), .B1(new_n934), .B2(new_n946), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n368), .C1(new_n960), .C2(new_n720), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n942), .A2(new_n696), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n698), .A2(new_n891), .A3(new_n720), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n933), .B(new_n513), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n963), .A2(new_n720), .A3(new_n925), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n962), .B1(new_n967), .B2(G148gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n959), .B1(new_n961), .B2(new_n968), .ZN(G1345gat));
  OAI21_X1  g768(.A(new_n384), .B1(new_n952), .B2(new_n857), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n958), .A2(new_n382), .A3(new_n383), .A4(new_n696), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1346gat));
  AOI21_X1  g771(.A(new_n385), .B1(new_n958), .B2(new_n759), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n650), .B1(new_n406), .B2(new_n407), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n960), .B2(new_n974), .ZN(G1347gat));
  NOR2_X1   g774(.A1(new_n723), .A2(new_n589), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI211_X1 g776(.A(new_n604), .B(new_n977), .C1(new_n856), .C2(new_n882), .ZN(new_n978));
  AOI21_X1  g777(.A(G169gat), .B1(new_n978), .B2(new_n811), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n977), .A2(new_n738), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n883), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n263), .A2(new_n270), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1348gat));
  NAND3_X1  g782(.A1(new_n978), .A2(new_n271), .A3(new_n720), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n981), .A2(new_n720), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(new_n271), .ZN(G1349gat));
  NAND3_X1  g785(.A1(new_n883), .A2(new_n696), .A3(new_n980), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n696), .A2(new_n313), .A3(new_n317), .ZN(new_n988));
  AOI22_X1  g787(.A1(new_n987), .A2(G183gat), .B1(new_n978), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g789(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n991));
  AND2_X1   g790(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n990), .A2(new_n993), .ZN(G1350gat));
  NAND3_X1  g793(.A1(new_n978), .A2(new_n320), .A3(new_n759), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n759), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n997), .B2(G190gat), .ZN(new_n998));
  AOI211_X1 g797(.A(KEYINPUT61), .B(new_n293), .C1(new_n981), .C2(new_n759), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G1351gat));
  NOR2_X1   g799(.A1(new_n784), .A2(new_n977), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n963), .A2(new_n966), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n891), .A2(G197gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n898), .A2(new_n513), .A3(new_n1001), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1004), .A2(new_n755), .ZN(new_n1005));
  OAI22_X1  g804(.A1(new_n1002), .A2(new_n1003), .B1(new_n1005), .B2(G197gat), .ZN(new_n1006));
  INV_X1    g805(.A(new_n1006), .ZN(G1352gat));
  NOR3_X1   g806(.A1(new_n1004), .A2(G204gat), .A3(new_n815), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n963), .A2(new_n720), .A3(new_n966), .ZN(new_n1010));
  INV_X1    g809(.A(new_n1001), .ZN(new_n1011));
  OAI21_X1  g810(.A(KEYINPUT127), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(G204gat), .ZN(new_n1013));
  NOR3_X1   g812(.A1(new_n1010), .A2(KEYINPUT127), .A3(new_n1011), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(G1353gat));
  INV_X1    g814(.A(new_n1004), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1016), .A2(new_n327), .A3(new_n696), .ZN(new_n1017));
  NAND4_X1  g816(.A1(new_n963), .A2(new_n696), .A3(new_n1001), .A4(new_n966), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(G1354gat));
  OAI21_X1  g821(.A(G218gat), .B1(new_n1002), .B2(new_n650), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1016), .A2(new_n328), .A3(new_n759), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(G1355gat));
endmodule


