//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT77), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT22), .B(G137), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT73), .ZN(new_n195));
  XNOR2_X1  g009(.A(G125), .B(G140), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(KEYINPUT16), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G125), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G140), .ZN(new_n201));
  AND4_X1   g015(.A1(new_n195), .A2(new_n199), .A3(new_n201), .A4(KEYINPUT16), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n197), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT74), .B1(new_n199), .B2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n198), .A4(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n204), .A3(G146), .A4(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(new_n201), .A3(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT73), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n199), .A2(new_n201), .A3(new_n195), .A4(KEYINPUT16), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n209), .A2(new_n212), .A3(G146), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n210), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G128), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT24), .B(G110), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT71), .B1(new_n222), .B2(G128), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT71), .B(new_n229), .C1(new_n222), .C2(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n223), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G110), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT72), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT72), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n234), .A3(G110), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n226), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n219), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G110), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n228), .A2(new_n238), .A3(new_n223), .A4(new_n230), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n224), .A2(new_n225), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n217), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT64), .A2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n196), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n214), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT76), .B1(new_n237), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n249));
  AOI211_X1 g063(.A(new_n249), .B(new_n246), .C1(new_n219), .C2(new_n236), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n194), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n219), .B2(new_n236), .ZN(new_n252));
  OR2_X1    g066(.A1(new_n252), .A2(new_n194), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT25), .B1(new_n254), .B2(new_n188), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n256), .B(G902), .C1(new_n251), .C2(new_n253), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n189), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT78), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(new_n189), .C1(new_n255), .C2(new_n257), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n189), .A2(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G122), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n268), .A2(KEYINPUT3), .A3(G107), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT79), .A2(G104), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT79), .A2(G104), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(G107), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(G107), .B1(new_n271), .B2(new_n272), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n270), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G101), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n222), .A2(G116), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G119), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT2), .B(G113), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n283), .A2(new_n284), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n283), .A2(new_n284), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT65), .A3(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n278), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n292));
  INV_X1    g106(.A(G101), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n273), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT80), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G107), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT79), .A2(G104), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT79), .A2(G104), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n269), .B1(new_n299), .B2(KEYINPUT3), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT80), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  AOI21_X1  g116(.A(G101), .B1(new_n302), .B2(G107), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n277), .B1(new_n276), .B2(G101), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n291), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n268), .A2(G107), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n293), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT5), .ZN(new_n310));
  OAI21_X1  g124(.A(G113), .B1(new_n280), .B2(KEYINPUT5), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n289), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g126(.A(new_n309), .B(new_n312), .C1(new_n295), .C2(new_n304), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n267), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n309), .B1(new_n295), .B2(new_n304), .ZN(new_n315));
  INV_X1    g129(.A(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n301), .B1(new_n300), .B2(new_n303), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n306), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n317), .B(new_n266), .C1(new_n321), .C2(new_n291), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n314), .A2(KEYINPUT6), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n243), .A2(G143), .A3(new_n244), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT0), .A2(G128), .ZN(new_n325));
  INV_X1    g139(.A(G143), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G146), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n326), .A2(G146), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT64), .B(G146), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT0), .B(G128), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G125), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n327), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n220), .B1(new_n324), .B2(KEYINPUT1), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n200), .B(new_n336), .C1(new_n337), .C2(new_n331), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n190), .A2(G224), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT82), .Z(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(new_n267), .C1(new_n307), .C2(new_n313), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n323), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n266), .B(KEYINPUT8), .Z(new_n346));
  INV_X1    g160(.A(new_n309), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n318), .B2(new_n319), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n312), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(new_n317), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n339), .B(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT83), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n346), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n315), .A2(new_n316), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n313), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n357));
  INV_X1    g171(.A(new_n351), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n339), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n360), .A3(new_n322), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n345), .A2(new_n361), .A3(new_n188), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n345), .A2(new_n361), .A3(new_n188), .A4(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G237), .A2(G953), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G214), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n326), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(G143), .A3(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT18), .A3(G131), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n245), .B1(new_n217), .B2(new_n196), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT18), .A2(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(KEYINPUT17), .A3(G131), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(G131), .ZN(new_n381));
  INV_X1    g195(.A(G131), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n372), .A2(new_n382), .A3(new_n373), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n384), .B2(KEYINPUT17), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n379), .B1(new_n219), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(new_n268), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n388), .B(new_n379), .C1(new_n219), .C2(new_n385), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT84), .A3(new_n188), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G475), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n390), .B2(new_n391), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT84), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n196), .B(KEYINPUT19), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n384), .B(new_n214), .C1(new_n398), .C2(new_n330), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n379), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n389), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n391), .ZN(new_n402));
  NOR2_X1   g216(.A1(G475), .A2(G902), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n404), .A2(KEYINPUT20), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(KEYINPUT20), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n394), .A2(new_n396), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(G234), .A2(G237), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n409), .A2(G952), .A3(new_n190), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT21), .B(G898), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT87), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n409), .A2(G902), .A3(G953), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n326), .A2(G128), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT13), .ZN(new_n418));
  OAI21_X1  g232(.A(KEYINPUT85), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT85), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n420), .A2(new_n326), .A3(KEYINPUT13), .A4(G128), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n220), .A2(G143), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n419), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G134), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n281), .A2(G122), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n281), .A2(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n296), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(G107), .ZN(new_n430));
  INV_X1    g244(.A(G134), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n423), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n425), .A2(new_n429), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n417), .B2(new_n423), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT86), .A3(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  INV_X1    g251(.A(new_n432), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n438), .B2(new_n434), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n426), .B(new_n427), .C1(KEYINPUT14), .C2(new_n296), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n428), .A2(new_n441), .A3(G107), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n439), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT9), .B(G234), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n446), .A2(new_n187), .A3(G953), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n444), .A2(new_n447), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n449), .A2(new_n450), .A3(G902), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n408), .A2(new_n416), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n369), .A2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n457));
  AND2_X1   g271(.A1(KEYINPUT64), .A2(G146), .ZN(new_n458));
  NOR2_X1   g272(.A1(KEYINPUT64), .A2(G146), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n326), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n329), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n332), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT66), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n431), .B2(G137), .ZN(new_n465));
  INV_X1    g279(.A(G137), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(KEYINPUT11), .A3(G134), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n431), .A2(G137), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G131), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n465), .A2(new_n467), .A3(new_n382), .A4(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT66), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n328), .B(new_n473), .C1(new_n331), .C2(new_n332), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n336), .B1(new_n337), .B2(new_n331), .ZN(new_n476));
  INV_X1    g290(.A(new_n468), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n431), .A2(G137), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n288), .A2(new_n290), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n370), .A2(G210), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT27), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G101), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(KEYINPUT29), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n475), .A2(new_n481), .ZN(new_n496));
  INV_X1    g310(.A(new_n482), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n483), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n499), .B2(KEYINPUT28), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n482), .B1(new_n475), .B2(new_n481), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n495), .B(KEYINPUT28), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n489), .B(new_n494), .C1(new_n500), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT28), .B1(new_n501), .B2(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n510), .A2(KEYINPUT70), .A3(new_n489), .A4(new_n494), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n476), .A2(new_n480), .ZN(new_n513));
  INV_X1    g327(.A(new_n472), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(new_n333), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n481), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n497), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n483), .ZN(new_n519));
  INV_X1    g333(.A(new_n493), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT29), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(new_n514), .A2(new_n333), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n482), .B1(new_n522), .B2(new_n481), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT28), .B1(new_n501), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n488), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n493), .B(KEYINPUT67), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n486), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n507), .A2(new_n511), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G472), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n518), .A2(new_n483), .A3(new_n493), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n518), .A2(KEYINPUT31), .A3(new_n483), .A4(new_n493), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n525), .A3(new_n486), .ZN(new_n535));
  INV_X1    g349(.A(new_n526), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT32), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n533), .A2(new_n534), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n536), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n538), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n530), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G110), .B(G140), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n190), .A2(G227), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n463), .A2(new_n278), .A3(new_n474), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n320), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n324), .A2(new_n327), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n220), .B1(new_n461), .B2(KEYINPUT1), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n336), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n347), .B(new_n555), .C1(new_n318), .C2(new_n319), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n476), .A2(KEYINPUT10), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n315), .A2(new_n559), .ZN(new_n560));
  AND4_X1   g374(.A1(new_n514), .A2(new_n552), .A3(new_n558), .A4(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n551), .A2(new_n320), .B1(new_n315), .B2(new_n559), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n514), .B1(new_n562), .B2(new_n558), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n550), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n556), .B1(new_n315), .B2(new_n476), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n472), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT12), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n514), .A3(new_n558), .ZN(new_n568));
  INV_X1    g382(.A(new_n550), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n570), .A3(new_n472), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n188), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n188), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n561), .A2(new_n563), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n569), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n567), .A2(new_n568), .A3(new_n571), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n550), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n575), .B(new_n577), .C1(new_n574), .C2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G221), .B1(new_n446), .B2(G902), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n265), .A2(new_n456), .A3(new_n547), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n584), .ZN(new_n588));
  OAI21_X1  g402(.A(G472), .B1(new_n537), .B2(G902), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n539), .B2(new_n537), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n265), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n362), .A2(new_n594), .A3(new_n364), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(new_n368), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n444), .A2(KEYINPUT90), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n447), .B1(new_n597), .B2(KEYINPUT91), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT90), .B1(new_n447), .B2(KEYINPUT91), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n445), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT33), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n452), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT89), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n444), .B(new_n448), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR4_X1   g420(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT89), .A4(KEYINPUT33), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n601), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT92), .B(G478), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT93), .B1(new_n451), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n604), .A2(new_n188), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  INV_X1    g426(.A(new_n609), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n407), .A2(new_n616), .A3(new_n416), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n365), .A2(KEYINPUT88), .A3(new_n366), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n596), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n596), .A2(new_n617), .A3(KEYINPUT94), .A4(new_n618), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n593), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND2_X1  g440(.A1(new_n596), .A2(new_n618), .ZN(new_n627));
  INV_X1    g441(.A(new_n454), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n408), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n593), .A2(new_n416), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n248), .A2(new_n250), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n262), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n259), .A2(new_n261), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n591), .A2(new_n456), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  AOI22_X1  g455(.A1(G472), .A2(new_n529), .B1(new_n540), .B2(new_n545), .ZN(new_n642));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n414), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n410), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n630), .A2(new_n585), .A3(new_n638), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n646), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n585), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n367), .B(KEYINPUT38), .ZN(new_n655));
  INV_X1    g469(.A(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n536), .A2(new_n499), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n531), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n546), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n407), .A2(new_n628), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n655), .A2(new_n368), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n638), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT95), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NOR2_X1   g479(.A1(new_n627), .A2(new_n642), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n407), .A2(new_n616), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n647), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n666), .A2(new_n585), .A3(new_n638), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  AOI21_X1  g484(.A(G902), .B1(new_n564), .B2(new_n572), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(new_n574), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n584), .A3(new_n575), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n264), .A2(new_n642), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n623), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NOR3_X1   g491(.A1(new_n627), .A2(new_n415), .A3(new_n629), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G116), .ZN(G18));
  AND2_X1   g494(.A1(new_n596), .A2(new_n618), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n673), .A2(new_n455), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n547), .A4(new_n638), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G119), .ZN(G21));
  NAND2_X1  g498(.A1(new_n264), .A2(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT96), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n259), .A2(new_n686), .A3(new_n261), .A4(new_n263), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n596), .A2(new_n618), .A3(new_n660), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n415), .A3(new_n673), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n526), .B1(new_n510), .B2(new_n489), .ZN(new_n691));
  INV_X1    g505(.A(new_n541), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n538), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n589), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n688), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NOR2_X1   g510(.A1(new_n627), .A2(new_n673), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n638), .A3(new_n668), .A4(new_n694), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  AOI21_X1  g513(.A(new_n642), .B1(new_n685), .B2(new_n687), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT97), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n580), .A2(new_n702), .A3(new_n550), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n579), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n580), .B2(new_n550), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n574), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n575), .A2(new_n577), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n584), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n365), .A2(new_n368), .A3(new_n366), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n701), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n584), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n581), .A2(KEYINPUT97), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(G469), .A3(new_n579), .A4(new_n703), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n576), .B1(new_n671), .B2(new_n574), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n365), .A2(new_n368), .A3(new_n366), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT98), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n668), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT99), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n264), .A2(new_n642), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n720), .A3(new_n721), .A4(new_n668), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n547), .A2(new_n261), .A3(new_n259), .A4(new_n263), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n710), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n720), .B1(new_n726), .B2(new_n668), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n719), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NOR2_X1   g543(.A1(new_n629), .A2(new_n647), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n715), .A2(KEYINPUT98), .A3(new_n716), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT98), .B1(new_n715), .B2(new_n716), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n721), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT100), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n718), .A2(new_n735), .A3(new_n721), .A4(new_n730), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n574), .B1(new_n582), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n579), .A4(new_n703), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n577), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n575), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT101), .ZN(new_n746));
  INV_X1    g560(.A(new_n743), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(KEYINPUT46), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n745), .A2(KEYINPUT101), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n584), .B(new_n651), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n408), .A2(new_n616), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT103), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT43), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n590), .A3(new_n638), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n709), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n752), .B(new_n761), .C1(new_n760), .C2(new_n759), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT105), .B(G137), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G39));
  NOR2_X1   g578(.A1(new_n748), .A2(new_n749), .ZN(new_n765));
  AND2_X1   g579(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n765), .A2(new_n711), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n765), .A2(new_n711), .B1(new_n768), .B2(new_n766), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n642), .A2(new_n264), .A3(new_n668), .A4(new_n716), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NAND2_X1  g586(.A1(new_n672), .A2(new_n575), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(KEYINPUT49), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n584), .A2(new_n368), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n753), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n655), .A2(new_n659), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n688), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n669), .A2(new_n698), .A3(new_n649), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n646), .B(KEYINPUT108), .Z(new_n782));
  NAND4_X1  g596(.A1(new_n259), .A2(new_n261), .A3(new_n637), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n689), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n659), .A3(new_n788), .A4(new_n715), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(new_n781), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n669), .A2(new_n698), .A3(new_n649), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n659), .A3(new_n715), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n786), .B2(new_n785), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n709), .A2(new_n628), .A3(new_n407), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n648), .A2(new_n585), .A3(new_n638), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n731), .A2(new_n732), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n638), .A2(new_n668), .A3(new_n694), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n735), .B1(new_n726), .B2(new_n730), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n733), .A2(KEYINPUT100), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n586), .A2(new_n683), .A3(new_n639), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n674), .B1(new_n623), .B2(new_n678), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n369), .B1(new_n667), .B2(new_n629), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n265), .A3(new_n591), .A4(new_n416), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n695), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT107), .B1(new_n812), .B2(new_n728), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n695), .A2(new_n586), .A3(new_n639), .A4(new_n683), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n675), .A2(new_n679), .A3(new_n810), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n802), .B1(new_n734), .B2(new_n736), .ZN(new_n817));
  AND4_X1   g631(.A1(KEYINPUT107), .A2(new_n728), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n797), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n820));
  OAI21_X1  g634(.A(new_n780), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n822));
  INV_X1    g636(.A(new_n815), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n586), .A2(new_n683), .A3(new_n639), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n688), .A2(new_n694), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n825), .B2(new_n690), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n817), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n719), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n722), .A2(new_n723), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n726), .A2(new_n668), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT99), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n822), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n728), .A2(new_n816), .A3(KEYINPUT107), .A4(new_n817), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n796), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n820), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT112), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n791), .B2(new_n793), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n790), .B2(new_n795), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n839), .A2(new_n794), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n833), .A2(new_n834), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n821), .B(new_n837), .C1(KEYINPUT53), .C2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n841), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n827), .A2(new_n832), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n845), .B(new_n849), .C1(new_n835), .C2(new_n836), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n756), .A2(new_n645), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n673), .A2(new_n709), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n638), .A2(new_n694), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n659), .A2(new_n645), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n265), .A3(new_n853), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n408), .A3(new_n615), .A4(new_n608), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n852), .A2(new_n825), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n655), .A2(new_n368), .A3(new_n673), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT50), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n767), .A2(new_n769), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n672), .A2(new_n711), .A3(new_n575), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n716), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n868), .B(KEYINPUT51), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n866), .B(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n859), .A3(new_n862), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n852), .A2(new_n700), .A3(new_n853), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(KEYINPUT48), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n861), .A2(new_n407), .A3(new_n616), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G952), .A3(new_n190), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n864), .B2(new_n697), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT48), .ZN(new_n890));
  INV_X1    g704(.A(new_n884), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT115), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(KEYINPUT115), .A2(new_n892), .A3(new_n885), .A4(new_n888), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n873), .B(new_n879), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n844), .A2(new_n851), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n779), .B1(new_n896), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n190), .A2(G952), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n323), .A2(new_n344), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT116), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n342), .B(KEYINPUT55), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n819), .A2(new_n820), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n188), .B1(new_n904), .B2(new_n849), .ZN(new_n905));
  AOI211_X1 g719(.A(KEYINPUT56), .B(new_n903), .C1(new_n905), .C2(G210), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n849), .B1(new_n835), .B2(new_n836), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(G210), .A3(G902), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n908), .B2(KEYINPUT117), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(KEYINPUT117), .B2(new_n908), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n899), .B(new_n906), .C1(new_n910), .C2(new_n903), .ZN(G51));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n188), .B(new_n742), .C1(new_n904), .C2(new_n849), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n576), .B(KEYINPUT118), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT57), .Z(new_n915));
  AOI21_X1  g729(.A(new_n845), .B1(new_n904), .B2(new_n849), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n851), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n573), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n918), .B2(new_n899), .ZN(new_n919));
  INV_X1    g733(.A(new_n899), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n850), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n922), .A2(new_n915), .B1(new_n564), .B2(new_n572), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT119), .B(new_n920), .C1(new_n923), .C2(new_n913), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G54));
  NAND2_X1  g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT120), .Z(new_n927));
  AND3_X1   g741(.A1(new_n905), .A2(new_n402), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n402), .B1(new_n905), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n899), .ZN(G60));
  OR2_X1    g744(.A1(new_n607), .A2(new_n606), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT59), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n922), .A2(new_n601), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n920), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n844), .B2(new_n851), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n931), .A2(new_n601), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n907), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n254), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n899), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(KEYINPUT61), .B1(new_n943), .B2(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n907), .A2(new_n636), .A3(new_n940), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G66));
  INV_X1    g761(.A(G224), .ZN(new_n948));
  OAI21_X1  g762(.A(G953), .B1(new_n413), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n811), .B(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n901), .B1(G898), .B2(new_n190), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  XNOR2_X1  g768(.A(new_n781), .B(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n664), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n629), .A2(new_n667), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n652), .A2(new_n960), .A3(new_n961), .A4(new_n709), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n721), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n771), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n958), .A2(new_n762), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n190), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n516), .A2(new_n517), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n398), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n700), .A2(new_n788), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n752), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n955), .A2(new_n737), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n762), .A2(new_n728), .A3(new_n771), .A4(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n976), .A2(new_n978), .A3(G953), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n969), .B1(G900), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n971), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G72));
  NOR2_X1   g798(.A1(new_n519), .A2(new_n493), .ZN(new_n985));
  INV_X1    g799(.A(new_n951), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n976), .A2(new_n978), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n965), .B2(new_n986), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n520), .B1(new_n518), .B2(new_n483), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(new_n994), .A3(new_n920), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n519), .A2(new_n520), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n990), .B1(new_n996), .B2(new_n531), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n995), .B1(new_n843), .B2(new_n997), .ZN(G57));
endmodule


