//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT2), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(KEYINPUT22), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G211gat), .B(G218gat), .Z(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT29), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n218), .A2(KEYINPUT79), .A3(KEYINPUT29), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n208), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n206), .B(new_n207), .Z(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n209), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n218), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n223), .A2(new_n228), .B1(G228gat), .B2(G233gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n208), .B1(new_n219), .B2(KEYINPUT3), .ZN(new_n230));
  AND4_X1   g029(.A1(G228gat), .A2(new_n228), .A3(G233gat), .A4(new_n230), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n229), .A2(new_n231), .A3(G22gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT80), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT80), .ZN(new_n234));
  XNOR2_X1  g033(.A(G78gat), .B(G106gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT31), .B(G50gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n229), .A2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G22gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n233), .A2(new_n234), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n237), .B(KEYINPUT78), .ZN(new_n241));
  INV_X1    g040(.A(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n232), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(G71gat), .ZN(new_n245));
  INV_X1    g044(.A(G99gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(G15gat), .B(G43gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT66), .B(G190gat), .Z(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT28), .ZN(new_n253));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT26), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n256), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n253), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n256), .A2(KEYINPUT23), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n256), .A2(KEYINPUT23), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(new_n262), .A3(new_n255), .ZN(new_n263));
  INV_X1    g062(.A(G183gat), .ZN(new_n264));
  INV_X1    g063(.A(G190gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT24), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT24), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(G183gat), .A3(G190gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(KEYINPUT25), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n264), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n250), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n280), .B2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n260), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n285), .A2(new_n286), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(G134gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n292), .B(new_n295), .C1(KEYINPUT1), .C2(new_n285), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n260), .ZN(new_n299));
  INV_X1    g098(.A(new_n283), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n281), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n291), .A2(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G227gat), .A2(G233gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n304), .B(KEYINPUT64), .Z(new_n305));
  NAND3_X1  g104(.A1(new_n298), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n249), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(KEYINPUT32), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n306), .B(KEYINPUT32), .C1(new_n307), .C2(new_n249), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n305), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n301), .A2(new_n302), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT34), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT34), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n310), .A3(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT35), .ZN(new_n325));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n302), .B1(KEYINPUT3), .B2(new_n208), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n225), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n302), .A2(new_n224), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT4), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n297), .A2(new_n208), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n329), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n297), .A2(new_n208), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(new_n327), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT0), .ZN(new_n345));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n334), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n339), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n343), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT6), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n343), .B2(new_n350), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT6), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n244), .A2(new_n324), .A3(new_n325), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n301), .A2(new_n226), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT73), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n284), .B2(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(new_n361), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n218), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n284), .A2(new_n363), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n301), .B2(new_n226), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n371), .A2(new_n372), .A3(new_n218), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(G64gat), .B(G92gat), .ZN(new_n377));
  XOR2_X1   g176(.A(new_n376), .B(new_n377), .Z(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n373), .B1(new_n218), .B2(new_n369), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n378), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT30), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n375), .A2(KEYINPUT30), .A3(new_n379), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n359), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n355), .B1(new_n353), .B2(KEYINPUT76), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n357), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n240), .A2(new_n243), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n312), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n324), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n312), .A2(new_n394), .A3(new_n320), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n384), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n386), .B1(new_n401), .B2(KEYINPUT35), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n356), .A2(new_n382), .A3(new_n357), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n218), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n364), .A2(new_n366), .A3(new_n406), .A4(new_n368), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(KEYINPUT84), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT37), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n218), .B1(new_n371), .B2(new_n372), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT38), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT85), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n381), .B2(new_n409), .ZN(new_n416));
  AND4_X1   g215(.A1(new_n415), .A2(new_n370), .A3(new_n374), .A4(new_n409), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n379), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n405), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT38), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT85), .B1(new_n375), .B2(KEYINPUT37), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n381), .A2(new_n415), .A3(new_n409), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n378), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n381), .A2(new_n409), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n330), .A2(new_n326), .A3(new_n340), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n328), .A2(new_n225), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n326), .B1(new_n349), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT39), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT81), .B(KEYINPUT39), .Z(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n347), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT40), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n437), .B1(new_n433), .B2(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n437), .C1(new_n433), .C2(new_n436), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n354), .B(new_n438), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n384), .A3(new_n383), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n244), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n403), .B1(new_n427), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n393), .B1(new_n385), .B2(new_n443), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(KEYINPUT86), .C1(new_n426), .C2(new_n419), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n399), .A2(KEYINPUT77), .A3(new_n390), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT77), .B1(new_n399), .B2(new_n390), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n393), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n322), .A2(new_n323), .B1(new_n394), .B2(new_n312), .ZN(new_n453));
  INV_X1    g252(.A(new_n397), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT36), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(KEYINPUT36), .B2(new_n324), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n402), .B1(new_n449), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G197gat), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT11), .B(G169gat), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n462), .B(KEYINPUT12), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT14), .ZN(new_n465));
  INV_X1    g264(.A(G29gat), .ZN(new_n466));
  INV_X1    g265(.A(G36gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G50gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G43gat), .ZN(new_n472));
  INV_X1    g271(.A(G43gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G50gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT15), .ZN(new_n475));
  NAND2_X1  g274(.A1(G29gat), .A2(G36gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n474), .A2(new_n478), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(KEYINPUT87), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n484), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n485), .A3(new_n469), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n475), .B1(new_n486), .B2(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n464), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n479), .B(new_n489), .C1(new_n478), .C2(new_n474), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n475), .A2(new_n476), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n470), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n486), .A2(new_n476), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(KEYINPUT89), .C1(new_n493), .C2(new_n475), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT16), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(G1gat), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G1gat), .B2(new_n496), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n495), .A2(new_n501), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT13), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n482), .A2(new_n487), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n501), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n511));
  NAND3_X1  g310(.A1(new_n488), .A2(new_n494), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT91), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n488), .A2(new_n494), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n505), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n516), .A2(new_n517), .A3(new_n503), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n507), .B1(new_n518), .B2(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  INV_X1    g319(.A(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n503), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n505), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n463), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n518), .A2(KEYINPUT18), .ZN(new_n529));
  INV_X1    g328(.A(new_n463), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n507), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(KEYINPUT92), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(new_n463), .C1(new_n519), .C2(new_n526), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT93), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n534), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n458), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G120gat), .B(G148gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT103), .ZN(new_n541));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  INV_X1    g344(.A(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G64gat), .ZN(new_n547));
  INV_X1    g346(.A(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G57gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n554), .B2(new_n550), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n545), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n554), .ZN(new_n558));
  INV_X1    g357(.A(G71gat), .ZN(new_n559));
  INV_X1    g358(.A(G78gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n561), .A2(new_n552), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT94), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT98), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(G85gat), .A3(G92gat), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n572), .A2(new_n574), .A3(KEYINPUT7), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT8), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n570), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n572), .A2(new_n574), .A3(KEYINPUT7), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n585), .A2(new_n569), .A3(new_n577), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n567), .A2(new_n568), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n557), .A3(new_n565), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n584), .A2(new_n563), .A3(new_n564), .A4(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n555), .A2(new_n556), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(KEYINPUT99), .A3(new_n587), .A4(new_n584), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n591), .B(KEYINPUT10), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n588), .A2(new_n557), .A3(new_n565), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n593), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT100), .B1(new_n601), .B2(new_n568), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n590), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n597), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n594), .A2(new_n593), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n592), .ZN(new_n608));
  INV_X1    g407(.A(new_n604), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n544), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n591), .B1(new_n608), .B2(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n568), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n589), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n604), .B1(new_n615), .B2(KEYINPUT101), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  AOI211_X1 g416(.A(new_n617), .B(new_n589), .C1(new_n613), .C2(new_n614), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT102), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n609), .B1(new_n603), .B2(new_n617), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(KEYINPUT101), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n610), .A2(new_n544), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT104), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n628), .B(new_n625), .C1(new_n619), .C2(new_n623), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n612), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n520), .A2(new_n509), .A3(new_n588), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n495), .B2(new_n588), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT97), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n631), .A2(new_n636), .A3(new_n634), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n638), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n638), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT21), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n501), .B1(new_n567), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n567), .A2(new_n648), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n653), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT95), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G183gat), .B(G211gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n657), .A2(new_n663), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n630), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n539), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n391), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n399), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n500), .B2(new_n673), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n675), .B(new_n676), .S(KEYINPUT42), .Z(G1325gat));
  OR2_X1    g476(.A1(new_n324), .A2(KEYINPUT36), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n455), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n670), .A2(G15gat), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(G15gat), .B1(new_n670), .B2(new_n324), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n244), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  INV_X1    g487(.A(new_n630), .ZN(new_n689));
  INV_X1    g488(.A(new_n666), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n647), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n539), .A2(new_n466), .A3(new_n391), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n458), .B2(new_n647), .ZN(new_n696));
  INV_X1    g495(.A(new_n647), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n452), .A2(new_n456), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n446), .B2(new_n448), .ZN(new_n699));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n697), .C1(new_n699), .C2(new_n402), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n532), .A2(new_n534), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n701), .A2(new_n391), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n694), .B1(new_n466), .B2(new_n704), .ZN(G1328gat));
  AOI211_X1 g504(.A(G36gat), .B(new_n399), .C1(KEYINPUT106), .C2(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n539), .A2(new_n692), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n701), .A2(new_n385), .A3(new_n703), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n467), .ZN(G1329gat));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n700), .A3(new_n679), .A4(new_n703), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G43gat), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT47), .B1(new_n713), .B2(KEYINPUT107), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n539), .A2(new_n692), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n324), .A2(new_n473), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n714), .B(new_n717), .ZN(G1330gat));
  NAND4_X1  g517(.A1(new_n701), .A2(G50gat), .A3(new_n393), .A4(new_n703), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n471), .B1(new_n715), .B2(new_n244), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g521(.A1(new_n449), .A2(new_n457), .ZN(new_n723));
  INV_X1    g522(.A(new_n402), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n702), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n689), .A2(new_n726), .A3(new_n667), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n390), .B(KEYINPUT108), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n546), .ZN(G1332gat));
  INV_X1    g531(.A(new_n728), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n399), .B(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n728), .B2(new_n456), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n324), .A2(new_n559), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1334gat));
  NOR2_X1   g548(.A1(new_n728), .A2(new_n244), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n560), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n726), .A2(new_n666), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n697), .B(new_n752), .C1(new_n699), .C2(new_n402), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n697), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n630), .A2(new_n580), .A3(new_n391), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT112), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n752), .A2(new_n630), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n701), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n391), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n763), .B2(new_n580), .ZN(G1336gat));
  NAND2_X1  g563(.A1(new_n735), .A2(new_n581), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n689), .B(new_n765), .C1(new_n755), .C2(new_n756), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n701), .A2(new_n735), .A3(new_n761), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n696), .A2(new_n700), .A3(new_n385), .A4(new_n761), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n771), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT113), .B1(new_n771), .B2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(new_n766), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(G1337gat));
  AOI21_X1  g575(.A(new_n689), .B1(new_n755), .B2(new_n756), .ZN(new_n777));
  AOI21_X1  g576(.A(G99gat), .B1(new_n777), .B2(new_n324), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n456), .A2(new_n246), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n762), .B2(new_n779), .ZN(G1338gat));
  XNOR2_X1  g579(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n244), .A2(G106gat), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n696), .A2(new_n700), .A3(new_n393), .A4(new_n761), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT114), .B(G106gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n783), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n784), .A2(KEYINPUT115), .A3(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(new_n782), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n689), .B(new_n792), .C1(new_n755), .C2(new_n756), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT115), .B1(new_n784), .B2(new_n787), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n668), .A2(new_n702), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT102), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n626), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n628), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n624), .A2(KEYINPUT104), .A3(new_n626), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n505), .B1(new_n522), .B2(new_n523), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n504), .A2(new_n506), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n462), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n531), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n645), .A2(new_n808), .A3(new_n646), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT54), .B1(new_n603), .B2(new_n604), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n619), .B2(new_n623), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n543), .B1(new_n605), .B2(KEYINPUT54), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT55), .B(new_n815), .C1(new_n816), .C2(new_n811), .ZN(new_n817));
  AND4_X1   g616(.A1(new_n804), .A2(new_n809), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n804), .A2(new_n726), .A3(new_n814), .A4(new_n817), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n630), .A2(new_n808), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n647), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n798), .B1(new_n822), .B2(new_n666), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT118), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n798), .C1(new_n822), .C2(new_n666), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n735), .A2(new_n390), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n244), .A2(new_n324), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n538), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n827), .A2(new_n730), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n398), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n735), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n702), .A2(G113gat), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT120), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n834), .A2(new_n840), .ZN(G1340gat));
  INV_X1    g640(.A(G120gat), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n831), .A2(new_n842), .A3(new_n689), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n837), .A2(new_n630), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n842), .ZN(G1341gat));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n294), .A3(new_n666), .ZN(new_n846));
  OAI21_X1  g645(.A(G127gat), .B1(new_n831), .B2(new_n690), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  OR3_X1    g647(.A1(new_n385), .A2(G134gat), .A3(new_n647), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n836), .A2(KEYINPUT56), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n831), .B2(new_n647), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT56), .B1(new_n836), .B2(new_n849), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n679), .A2(new_n244), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n538), .A2(G141gat), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n835), .A2(new_n736), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT121), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n829), .A2(new_n456), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n804), .A2(new_n814), .A3(new_n817), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n820), .B1(new_n860), .B2(new_n538), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n647), .ZN(new_n862));
  INV_X1    g661(.A(new_n818), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n666), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n798), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n393), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n859), .B1(new_n866), .B2(KEYINPUT57), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n824), .A2(new_n868), .A3(new_n393), .A4(new_n826), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n726), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n858), .B1(new_n870), .B2(G141gat), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n867), .A2(new_n869), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n538), .ZN(new_n874));
  INV_X1    g673(.A(new_n854), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n827), .A2(new_n730), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n736), .A4(new_n855), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n857), .A2(new_n871), .B1(new_n879), .B2(new_n858), .ZN(G1344gat));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n876), .A2(new_n881), .A3(new_n630), .A4(new_n736), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n393), .A2(new_n868), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n534), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n535), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n804), .A3(new_n814), .A4(new_n817), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n697), .B1(new_n887), .B2(new_n820), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n690), .B1(new_n888), .B2(new_n818), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n668), .A2(new_n538), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n829), .A2(new_n456), .A3(new_n630), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n824), .A2(new_n393), .A3(new_n826), .ZN(new_n895));
  AOI211_X1 g694(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n881), .B1(new_n896), .B2(KEYINPUT125), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n893), .B1(new_n895), .B2(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n894), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n883), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n630), .A3(new_n869), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n904), .B2(new_n906), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n882), .B1(new_n903), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n873), .B2(new_n690), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n876), .A2(new_n736), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n666), .A2(new_n203), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1346gat));
  OAI21_X1  g713(.A(G162gat), .B1(new_n873), .B2(new_n647), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n876), .A2(new_n204), .A3(new_n399), .A4(new_n697), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n729), .A2(new_n399), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n828), .A2(new_n830), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(G169gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n919), .A2(new_n920), .A3(new_n538), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n827), .A2(new_n391), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n398), .A3(new_n735), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n726), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n925), .B2(new_n920), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n919), .B2(new_n689), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n689), .A2(G176gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n923), .B2(new_n928), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n919), .B2(new_n690), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n666), .A2(new_n251), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n923), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n930), .B(new_n934), .C1(new_n923), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n919), .B2(new_n647), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT61), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n697), .A2(new_n250), .ZN(new_n940));
  OR3_X1    g739(.A1(new_n923), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n923), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n938), .A2(new_n943), .ZN(G1351gat));
  NOR2_X1   g743(.A1(new_n875), .A2(new_n736), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n824), .A2(new_n390), .A3(new_n945), .A4(new_n826), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n726), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n918), .A2(new_n456), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n893), .B(new_n949), .C1(new_n895), .C2(KEYINPUT57), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n886), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n898), .A2(new_n456), .A3(new_n918), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n953), .B2(new_n689), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n689), .A2(G204gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n946), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n954), .A2(new_n955), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n961), .B1(new_n950), .B2(new_n630), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n959), .A2(new_n958), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT127), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n960), .A2(new_n964), .ZN(G1353gat));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n211), .A3(new_n666), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n666), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n967), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n953), .B2(new_n647), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n947), .A2(new_n212), .A3(new_n697), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1355gat));
endmodule


