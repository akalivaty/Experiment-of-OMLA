//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G143), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT66), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n196), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT17), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT77), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT77), .A4(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n192), .A2(KEYINPUT17), .A3(new_n197), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G113), .B(G122), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT90), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT18), .A3(G131), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n191), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n191), .A2(new_n222), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(new_n206), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n210), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(new_n210), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n223), .B(new_n224), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n217), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n220), .B1(new_n217), .B2(new_n230), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n187), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT92), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT92), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n235), .B(new_n187), .C1(new_n231), .C2(new_n232), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(G475), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n198), .A2(new_n200), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n225), .B(KEYINPUT19), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n212), .B1(new_n239), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n230), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n220), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n217), .A2(new_n220), .A3(new_n230), .ZN(new_n244));
  AOI21_X1  g058(.A(G475), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT91), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n187), .B(new_n245), .C1(new_n246), .C2(KEYINPUT20), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(KEYINPUT20), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n187), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n237), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G122), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT14), .B1(new_n252), .B2(G116), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT14), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G122), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n253), .B(new_n256), .C1(new_n255), .C2(G122), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G107), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT97), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n255), .A2(G122), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n252), .A2(G116), .ZN(new_n261));
  OR3_X1    g075(.A1(new_n260), .A2(new_n261), .A3(G107), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(G134), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(G143), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(KEYINPUT96), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(KEYINPUT96), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n259), .A2(new_n262), .A3(new_n273), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT13), .B1(new_n265), .B2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n266), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT93), .B(new_n269), .C1(new_n264), .C2(KEYINPUT13), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n264), .A2(KEYINPUT13), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G107), .B1(new_n260), .B2(new_n261), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(G134), .B1(new_n282), .B2(new_n262), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n271), .B(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n283), .A2(KEYINPUT95), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT95), .B1(new_n283), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n275), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT9), .B(G234), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G217), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n290), .A2(new_n291), .A3(G953), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n275), .B(new_n292), .C1(new_n286), .C2(new_n287), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(KEYINPUT98), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n288), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT98), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n292), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n187), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G478), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n302), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n296), .A2(new_n299), .A3(new_n187), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n189), .A2(G952), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(G234), .B2(G237), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT21), .B(G898), .Z(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n187), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n251), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(new_n187), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n210), .B2(G143), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n210), .A2(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT1), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n210), .A3(G143), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n320), .A2(new_n321), .A3(G128), .A4(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n265), .A2(G146), .ZN(new_n324));
  OAI21_X1  g138(.A(G128), .B1(new_n324), .B2(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n265), .A2(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g145(.A(G107), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G104), .ZN(new_n333));
  INV_X1    g147(.A(G101), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n219), .A2(G107), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n332), .A2(G104), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n219), .A2(G107), .ZN(new_n338));
  OAI21_X1  g152(.A(G101), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n339), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT65), .B1(new_n265), .B2(G146), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n322), .B1(new_n343), .B2(new_n324), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n325), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n323), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT11), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n270), .B2(G137), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n270), .A2(G137), .ZN(new_n351));
  INV_X1    g165(.A(G137), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT11), .A3(G134), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G131), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n199), .A2(new_n351), .A3(new_n350), .A4(new_n353), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT67), .B1(new_n354), .B2(G131), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT12), .B1(new_n347), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n345), .A2(new_n323), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(new_n342), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n336), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n265), .A2(KEYINPUT65), .A3(G146), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n319), .B2(new_n318), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT0), .A2(G128), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(KEYINPUT64), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT0), .A2(G128), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n319), .B2(new_n326), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n368), .A2(new_n370), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(new_n375), .A3(G101), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n340), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n363), .A2(new_n359), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT12), .ZN(new_n380));
  OAI221_X1 g194(.A(new_n380), .B1(new_n357), .B2(new_n358), .C1(new_n341), .C2(new_n346), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n360), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  XOR2_X1   g196(.A(G110), .B(G140), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n189), .A2(G227), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n359), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(new_n378), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n346), .A2(KEYINPUT10), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n387), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n379), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(G469), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n392), .B2(new_n379), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n360), .A2(new_n379), .A3(new_n393), .A4(new_n381), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n398), .B(new_n187), .C1(new_n400), .C2(new_n396), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n316), .B(new_n395), .C1(new_n401), .C2(G469), .ZN(new_n402));
  OAI21_X1  g216(.A(G221), .B1(new_n290), .B2(G902), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G214), .B1(G237), .B2(G902), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT84), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n371), .A2(new_n373), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n320), .A2(new_n322), .A3(new_n370), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n408), .A2(G125), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(G125), .B1(new_n323), .B2(new_n328), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT7), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n374), .A2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n329), .A2(new_n205), .ZN(new_n414));
  INV_X1    g228(.A(G224), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n410), .B2(new_n411), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT7), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT88), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT87), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n255), .A2(KEYINPUT5), .A3(G119), .ZN(new_n423));
  INV_X1    g237(.A(G113), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G116), .B(G119), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT5), .ZN(new_n427));
  INV_X1    g241(.A(G119), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G116), .ZN(new_n429));
  OAI211_X1 g243(.A(KEYINPUT87), .B(G113), .C1(new_n429), .C2(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(KEYINPUT2), .A2(G113), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n255), .A2(G119), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT2), .A2(G113), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n432), .A2(new_n429), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n342), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n429), .A2(new_n433), .A3(KEYINPUT5), .ZN(new_n437));
  OAI21_X1  g251(.A(G113), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n340), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT8), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n421), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  NOR4_X1   g259(.A1(new_n436), .A2(new_n440), .A3(KEYINPUT88), .A4(new_n443), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n412), .B(new_n420), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT89), .ZN(new_n448));
  INV_X1    g262(.A(new_n436), .ZN(new_n449));
  INV_X1    g263(.A(new_n439), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n342), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n444), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT88), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n441), .A2(new_n421), .A3(new_n444), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n412), .A4(new_n420), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n432), .B(new_n434), .C1(new_n426), .C2(KEYINPUT69), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n432), .A2(new_n434), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n429), .A2(new_n433), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n366), .A2(new_n463), .A3(new_n376), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n450), .A2(new_n340), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(new_n465), .A3(new_n442), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n448), .A2(new_n457), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n418), .A2(new_n419), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n442), .B1(new_n464), .B2(new_n465), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(KEYINPUT86), .A3(new_n471), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n466), .A2(new_n470), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT85), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n479));
  NOR4_X1   g293(.A1(new_n466), .A2(new_n470), .A3(new_n479), .A4(new_n471), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n469), .B(new_n476), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n468), .A2(new_n481), .A3(new_n187), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n468), .A2(new_n481), .A3(new_n187), .A4(new_n483), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n407), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n313), .A2(new_n404), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n291), .B1(G234), .B2(new_n187), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n227), .A2(new_n212), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT73), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n263), .B2(G119), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n263), .A2(G119), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n428), .A2(KEYINPUT73), .A3(G128), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT74), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n495), .A2(new_n497), .A3(new_n500), .A4(new_n496), .ZN(new_n501));
  OR2_X1    g315(.A1(KEYINPUT24), .A2(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT24), .A2(G110), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(KEYINPUT75), .A3(new_n503), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n499), .A2(new_n501), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT76), .B1(new_n428), .B2(G128), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT23), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n428), .A2(G128), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n496), .A2(KEYINPUT76), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(G110), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n493), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n493), .B(KEYINPUT78), .C1(new_n508), .C2(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n499), .A2(new_n501), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n506), .A2(new_n507), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n514), .A2(G110), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n213), .A3(new_n214), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n522), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n514), .A2(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT78), .B1(new_n531), .B2(new_n493), .ZN(new_n532));
  INV_X1    g346(.A(new_n519), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT79), .B(new_n525), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT22), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G137), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n528), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT79), .B(new_n538), .C1(new_n520), .C2(new_n525), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT25), .B1(new_n542), .B2(new_n187), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT80), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n492), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n538), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT79), .B1(new_n520), .B2(new_n525), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n187), .B1(new_n548), .B2(new_n540), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT25), .B(new_n187), .C1(new_n548), .C2(new_n540), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n545), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n374), .B1(new_n357), .B2(new_n358), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n352), .A2(G134), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n270), .A2(G137), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n354), .B2(new_n197), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT68), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n356), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n329), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(KEYINPUT70), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n356), .A2(new_n568), .A3(new_n559), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n329), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n565), .B1(new_n556), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n463), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n463), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n556), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT27), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT26), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n334), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n572), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT31), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(KEYINPUT28), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT28), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n556), .A2(new_n570), .A3(new_n582), .A4(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n556), .A2(new_n564), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n463), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n577), .B(G101), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(KEYINPUT71), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT71), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n581), .A2(new_n583), .B1(new_n463), .B2(new_n585), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n572), .A2(new_n593), .A3(new_n578), .A4(new_n574), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n580), .A2(new_n589), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G472), .A2(G902), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(KEYINPUT32), .A3(new_n596), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n587), .A2(new_n588), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n578), .B1(new_n572), .B2(new_n574), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(KEYINPUT29), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n556), .A2(new_n570), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n584), .B1(new_n573), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n578), .A2(KEYINPUT29), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n187), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G472), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n599), .A2(new_n600), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n491), .A2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n542), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n555), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n313), .A2(KEYINPUT99), .A3(new_n404), .A4(new_n487), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n490), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  AND3_X1   g429(.A1(new_n555), .A2(new_n404), .A3(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n485), .A2(new_n486), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n405), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n296), .A2(new_n619), .A3(new_n299), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n294), .A2(KEYINPUT33), .A3(new_n295), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n294), .A2(KEYINPUT100), .A3(KEYINPUT33), .A4(new_n295), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n301), .A2(G902), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n620), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n300), .A2(new_n301), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n251), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n618), .A2(new_n312), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n595), .A2(new_n187), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n631), .A2(G472), .B1(new_n596), .B2(new_n595), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n616), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n405), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n636), .B(new_n312), .C1(new_n485), .C2(new_n486), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n234), .A2(new_n236), .ZN(new_n638));
  AOI22_X1  g452(.A1(G475), .A2(new_n638), .B1(new_n303), .B2(new_n305), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n249), .B(KEYINPUT20), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n616), .A3(new_n632), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n332), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT101), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT35), .ZN(G9));
  NOR2_X1   g459(.A1(new_n538), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n526), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n610), .ZN(new_n648));
  INV_X1    g462(.A(new_n492), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n549), .A2(new_n544), .A3(new_n550), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n649), .B(new_n650), .C1(new_n651), .C2(new_n543), .ZN(new_n652));
  INV_X1    g466(.A(new_n554), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n490), .A3(new_n613), .A4(new_n632), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT103), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AND2_X1   g476(.A1(new_n609), .A2(new_n404), .ZN(new_n663));
  INV_X1    g477(.A(new_n306), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT104), .B(G900), .Z(new_n665));
  AOI21_X1  g479(.A(new_n308), .B1(new_n311), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n640), .A2(new_n237), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n618), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT102), .B1(new_n555), .B2(new_n648), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n663), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XNOR2_X1  g487(.A(new_n666), .B(KEYINPUT39), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n404), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT107), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n654), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n604), .A2(new_n573), .ZN(new_n682));
  INV_X1    g496(.A(new_n574), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n588), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n579), .A2(G472), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(G472), .A2(G902), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT105), .Z(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n599), .A3(new_n600), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT106), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n617), .B(KEYINPUT38), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n251), .A2(new_n306), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n691), .A2(new_n405), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n680), .A2(new_n681), .A3(new_n690), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND3_X1  g509(.A1(new_n628), .A2(new_n251), .A3(new_n667), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT108), .B1(new_n618), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n250), .A2(new_n247), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n699), .A2(new_n237), .B1(new_n626), .B2(new_n627), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n636), .B1(new_n485), .B2(new_n486), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n667), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n663), .C1(new_n670), .C2(new_n671), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  OR2_X1    g520(.A1(new_n401), .A2(G469), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n401), .A2(G469), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n403), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n612), .A2(KEYINPUT109), .A3(new_n630), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n555), .A2(new_n609), .A3(new_n711), .A4(new_n611), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n637), .A2(new_n700), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT41), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G113), .ZN(G15));
  NAND3_X1  g533(.A1(new_n641), .A2(new_n612), .A3(new_n711), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  AND2_X1   g535(.A1(new_n711), .A2(new_n701), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n609), .A2(new_n313), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n658), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n605), .A2(new_n588), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n580), .A3(new_n594), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n631), .A2(G472), .B1(new_n596), .B2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n555), .A2(new_n611), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n711), .A2(new_n692), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n637), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n637), .A2(new_n555), .A3(new_n611), .A4(new_n728), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT110), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT111), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n252), .ZN(G24));
  INV_X1    g552(.A(new_n696), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n722), .A2(new_n654), .A3(new_n739), .A4(new_n728), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND3_X1  g555(.A1(new_n485), .A2(new_n486), .A3(new_n405), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n316), .B1(new_n401), .B2(G469), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n388), .B2(new_n394), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT112), .B1(new_n382), .B2(new_n387), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n314), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n403), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n612), .A2(KEYINPUT42), .A3(new_n739), .A4(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n555), .A3(new_n609), .A4(new_n611), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n696), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  INV_X1    g569(.A(new_n752), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n668), .A2(new_n664), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  INV_X1    g573(.A(new_n654), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n632), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n628), .A2(new_n237), .A3(new_n699), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT43), .Z(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n745), .A2(new_n746), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n314), .B1(new_n767), .B2(KEYINPUT45), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n388), .A2(new_n394), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n316), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n707), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n403), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n674), .ZN(new_n778));
  INV_X1    g592(.A(new_n742), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n761), .A2(new_n763), .A3(KEYINPUT44), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n766), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NAND2_X1  g596(.A1(new_n777), .A2(KEYINPUT47), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n555), .A2(new_n611), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n609), .A3(new_n696), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(new_n403), .C1(new_n775), .C2(new_n776), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n779), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(new_n690), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n784), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n709), .B(KEYINPUT113), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n797), .A2(new_n710), .A3(new_n691), .A4(new_n762), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n791), .A2(new_n796), .A3(new_n406), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n783), .A2(new_n787), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n403), .B2(new_n792), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n729), .A2(new_n308), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(new_n763), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n803), .A2(KEYINPUT117), .A3(new_n779), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n779), .A3(new_n763), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n711), .A2(new_n636), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n691), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n802), .A2(new_n812), .A3(new_n763), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT50), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n711), .A2(new_n779), .A3(new_n308), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n763), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT119), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n763), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n654), .A2(new_n728), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n821), .A2(new_n822), .B1(new_n814), .B2(KEYINPUT50), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n628), .A2(new_n251), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n791), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n808), .A2(new_n815), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT48), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n821), .B2(new_n612), .ZN(new_n830));
  INV_X1    g644(.A(new_n612), .ZN(new_n831));
  AOI211_X1 g645(.A(KEYINPUT48), .B(new_n831), .C1(new_n818), .C2(new_n820), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n803), .A2(new_n722), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n790), .A2(new_n784), .A3(new_n700), .A4(new_n816), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(G952), .A3(new_n189), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(KEYINPUT120), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n823), .A2(new_n825), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT51), .A3(new_n815), .A4(new_n808), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n836), .B(new_n834), .C1(new_n830), .C2(new_n832), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n828), .A2(new_n837), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(new_n654), .A2(new_n739), .A3(new_n728), .A4(new_n749), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n844), .A2(new_n845), .B1(new_n756), .B2(new_n757), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n654), .A2(new_n739), .A3(new_n728), .A4(new_n749), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n668), .A2(new_n306), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n658), .A2(new_n663), .A3(new_n779), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n659), .A2(new_n736), .A3(new_n717), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n639), .A2(new_n699), .B1(new_n628), .B2(new_n251), .ZN(new_n853));
  INV_X1    g667(.A(new_n487), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n853), .A2(new_n854), .A3(new_n312), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n616), .A3(new_n632), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(new_n614), .A3(new_n720), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n658), .A2(new_n722), .A3(new_n723), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n851), .A2(new_n852), .A3(new_n754), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n692), .A2(new_n617), .A3(new_n405), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n748), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n760), .A3(new_n667), .A4(new_n689), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n705), .A2(new_n672), .A3(new_n740), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT52), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n658), .B(new_n663), .C1(new_n669), .C2(new_n704), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n740), .A4(new_n864), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n860), .A2(new_n861), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n866), .A2(new_n869), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n846), .A2(new_n754), .A3(new_n850), .A4(new_n848), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n659), .A2(new_n736), .A3(new_n717), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n724), .A2(new_n614), .A3(new_n720), .A4(new_n856), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT54), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n861), .B1(new_n860), .B2(new_n870), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n876), .A3(KEYINPUT53), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n879), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n882), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n843), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n799), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT121), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n799), .C1(new_n887), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(G75));
  AOI21_X1  g707(.A(new_n187), .B1(new_n880), .B2(new_n882), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G210), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  INV_X1    g710(.A(new_n478), .ZN(new_n897));
  INV_X1    g711(.A(new_n480), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n897), .A2(new_n898), .B1(new_n474), .B2(new_n475), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(new_n469), .Z(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n895), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n189), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  AND2_X1   g719(.A1(new_n878), .A2(new_n883), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n315), .B(KEYINPUT57), .Z(new_n907));
  OAI221_X1 g721(.A(new_n398), .B1(new_n396), .B2(new_n400), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n894), .A2(new_n770), .A3(new_n768), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n243), .A2(new_n244), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n914), .A2(new_n915), .A3(new_n904), .ZN(G60));
  NAND3_X1  g730(.A1(new_n620), .A2(new_n624), .A3(new_n623), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  NOR3_X1   g733(.A1(new_n906), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n884), .A2(new_n886), .A3(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n904), .B(new_n920), .C1(new_n917), .C2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  AOI21_X1  g739(.A(new_n542), .B1(new_n885), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n904), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n885), .A2(new_n647), .A3(new_n925), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n927), .A2(new_n928), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n929));
  NOR2_X1   g743(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G66));
  OAI21_X1  g745(.A(G953), .B1(new_n310), .B2(new_n415), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n874), .A2(new_n875), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(G953), .ZN(new_n934));
  INV_X1    g748(.A(new_n899), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(G898), .B2(new_n189), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n934), .B(new_n936), .ZN(G69));
  NOR2_X1   g751(.A1(new_n566), .A2(new_n571), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n239), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OR4_X1    g754(.A1(new_n831), .A2(new_n677), .A3(new_n742), .A4(new_n853), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n781), .A2(new_n788), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n867), .A2(new_n740), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n694), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n694), .A2(new_n944), .A3(KEYINPUT62), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n940), .B1(new_n949), .B2(G953), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(KEYINPUT123), .B(new_n940), .C1(new_n949), .C2(G953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n766), .A2(new_n779), .A3(new_n780), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n831), .B2(new_n862), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n778), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n944), .A2(new_n788), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n754), .A2(new_n758), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n958), .A2(new_n189), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(G900), .A2(G953), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n939), .A3(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n952), .A2(new_n954), .A3(new_n955), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT124), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n961), .A2(KEYINPUT124), .A3(new_n939), .A4(new_n962), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n952), .A2(new_n966), .A3(new_n955), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n968), .A2(new_n969), .A3(new_n953), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n968), .B2(new_n953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(G72));
  NAND3_X1  g786(.A1(new_n572), .A2(new_n574), .A3(new_n588), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n958), .A2(new_n933), .A3(new_n959), .A4(new_n960), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n686), .B(KEYINPUT63), .Z(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n975), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n949), .B2(new_n933), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n572), .A2(new_n574), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n578), .ZN(new_n980));
  OAI22_X1  g794(.A1(new_n978), .A2(new_n980), .B1(G952), .B2(new_n189), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n885), .A2(new_n975), .A3(new_n973), .A4(new_n980), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n976), .B(new_n981), .C1(new_n984), .C2(new_n985), .ZN(G57));
endmodule


