//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G146), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT66), .B1(new_n188), .B2(G143), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n193), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n189), .A2(new_n190), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n193), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n198), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n207), .A2(G134), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT67), .A2(G131), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT67), .A2(G131), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n208), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT67), .A2(G131), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n205), .A2(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT67), .A2(G131), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  OR3_X1    g036(.A1(new_n205), .A2(KEYINPUT69), .A3(G137), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n205), .B2(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G131), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n203), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n206), .A2(new_n208), .A3(new_n218), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G131), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n188), .A2(G143), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT65), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT65), .A2(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n231), .B1(new_n234), .B2(G143), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT0), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(new_n196), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n196), .A3(KEYINPUT64), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n195), .A2(new_n194), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n191), .A3(new_n237), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n227), .A2(KEYINPUT70), .B1(new_n230), .B2(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n215), .A2(new_n221), .B1(G131), .B2(new_n225), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n203), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT30), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n251), .B2(G119), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n253));
  INV_X1    g067(.A(G119), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G116), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n252), .A2(new_n255), .B1(new_n251), .B2(G119), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT2), .B(G113), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n203), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(KEYINPUT72), .B(new_n198), .C1(new_n199), .C2(new_n202), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n260), .A2(new_n247), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n215), .A2(new_n221), .B1(G131), .B2(new_n228), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n242), .A2(new_n244), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT30), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n258), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n250), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G237), .ZN(new_n271));
  AOI21_X1  g085(.A(G953), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G210), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n272), .B2(G210), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT26), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n274), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n277), .A2(new_n280), .A3(G101), .ZN(new_n281));
  AOI21_X1  g095(.A(G101), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n260), .A2(new_n247), .A3(new_n261), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n230), .A2(new_n245), .ZN(new_n285));
  INV_X1    g099(.A(new_n258), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT74), .B1(new_n267), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n227), .A2(KEYINPUT70), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n249), .A3(new_n285), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n265), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n286), .B1(new_n294), .B2(new_n284), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n287), .ZN(new_n297));
  INV_X1    g111(.A(G101), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n279), .B1(new_n278), .B2(new_n274), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT26), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n277), .A2(new_n280), .A3(G101), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n296), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n288), .B1(new_n293), .B2(new_n295), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n291), .A2(new_n258), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n287), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n284), .A2(KEYINPUT28), .A3(new_n285), .A4(new_n286), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n308), .A2(new_n309), .B1(new_n314), .B2(new_n303), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G472), .A2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT32), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n317), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n307), .B2(new_n315), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n323), .B2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g138(.A(G472), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n310), .A2(new_n312), .A3(new_n283), .A4(new_n313), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n297), .B1(new_n293), .B2(new_n295), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n283), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n284), .A2(new_n285), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n258), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n312), .A2(new_n313), .A3(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n303), .A2(new_n327), .ZN(new_n333));
  AOI21_X1  g147(.A(G902), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n325), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n323), .B2(KEYINPUT32), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n321), .A2(new_n324), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n254), .B2(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(new_n340), .C1(G119), .C2(new_n196), .ZN(new_n341));
  XNOR2_X1  g155(.A(G119), .B(G128), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT24), .B(G110), .Z(new_n343));
  AOI22_X1  g157(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(new_n188), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n349), .A2(KEYINPUT16), .A3(G140), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G146), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n344), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n341), .A2(G110), .B1(new_n342), .B2(new_n343), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(G146), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n234), .A2(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G953), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(G221), .A3(G234), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n365), .A2(KEYINPUT22), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(KEYINPUT22), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n207), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n368), .B(G137), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n358), .A3(new_n362), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n370), .A2(KEYINPUT25), .A3(new_n371), .A4(new_n373), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT76), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G217), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(G234), .B2(new_n371), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT76), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n381), .A3(new_n375), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n370), .A2(new_n373), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT77), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n380), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n390));
  OAI21_X1  g204(.A(G128), .B1(new_n200), .B2(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n232), .A2(new_n233), .A3(new_n193), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n195), .A2(new_n194), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n198), .ZN(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G101), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT79), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n399), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n398), .A2(G104), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n396), .A2(G107), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n410), .A3(new_n298), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n395), .A2(new_n401), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n401), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n399), .A2(new_n406), .B1(new_n400), .B2(new_n405), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(new_n298), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n203), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n230), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT12), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n260), .A2(KEYINPUT10), .A3(new_n261), .A4(new_n415), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n196), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n243), .B2(new_n191), .ZN(new_n421));
  AND4_X1   g235(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n197), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n401), .B(new_n411), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n409), .B1(new_n403), .B2(new_n405), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n397), .A2(new_n399), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n426), .B(G101), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G101), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n411), .A3(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n245), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n419), .A2(new_n263), .A3(new_n425), .A4(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n364), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n411), .A2(new_n401), .ZN(new_n438));
  OAI21_X1  g252(.A(G128), .B1(new_n392), .B2(new_n390), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n235), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n440), .A3(new_n198), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n423), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT12), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n230), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n418), .A2(new_n433), .A3(new_n437), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n443), .B1(new_n442), .B2(new_n230), .ZN(new_n447));
  AOI211_X1 g261(.A(KEYINPUT12), .B(new_n263), .C1(new_n441), .C2(new_n423), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n433), .A4(new_n437), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT10), .B1(new_n415), .B2(new_n395), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n431), .A2(new_n429), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(new_n245), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n263), .B1(new_n454), .B2(new_n419), .ZN(new_n455));
  INV_X1    g269(.A(new_n433), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n436), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT80), .B(G469), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n371), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n437), .B1(new_n455), .B2(new_n456), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n449), .A2(new_n433), .A3(new_n436), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n371), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G469), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT9), .B(G234), .ZN(new_n467));
  OAI21_X1  g281(.A(G221), .B1(new_n467), .B2(G902), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT78), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G214), .B1(G237), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n349), .B(new_n198), .C1(new_n199), .C2(new_n202), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n349), .B1(new_n242), .B2(new_n244), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT84), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n476), .A2(KEYINPUT84), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G224), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n431), .A2(new_n258), .A3(new_n429), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n256), .ZN(new_n489));
  INV_X1    g303(.A(G113), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n251), .A2(G119), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n489), .A2(new_n492), .B1(new_n257), .B2(new_n256), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n415), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G122), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n486), .A2(new_n494), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n495), .A2(KEYINPUT83), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n496), .A2(KEYINPUT6), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n497), .A2(KEYINPUT6), .A3(new_n498), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n485), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n256), .A2(new_n257), .ZN(new_n502));
  INV_X1    g316(.A(new_n492), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n415), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n493), .A2(new_n438), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n495), .B(KEYINPUT8), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n483), .A2(KEYINPUT7), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n475), .B2(new_n476), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n509), .A2(new_n496), .A3(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT7), .A4(new_n483), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(new_n514), .A3(new_n516), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n473), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n471), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n270), .A2(G237), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n525));
  OAI211_X1 g339(.A(G214), .B(new_n364), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(new_n193), .ZN(new_n527));
  AOI21_X1  g341(.A(G143), .B1(new_n272), .B2(G214), .ZN(new_n528));
  NAND2_X1  g342(.A1(KEYINPUT18), .A2(G131), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT86), .Z(new_n530));
  OR3_X1    g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n361), .B1(new_n188), .B2(new_n355), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n193), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n272), .A2(G143), .A3(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n529), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(KEYINPUT85), .B(new_n529), .C1(new_n534), .C2(new_n535), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n531), .B(new_n532), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT87), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n396), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n352), .A2(new_n188), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n360), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n211), .A2(new_n212), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n534), .B2(new_n535), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(KEYINPUT17), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n546), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n527), .B2(new_n528), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n534), .A2(new_n546), .A3(new_n535), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n540), .A2(new_n543), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n552), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n355), .B(KEYINPUT19), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n234), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n360), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n543), .B1(new_n540), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n523), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(G475), .A2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n543), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n532), .B1(new_n536), .B2(new_n530), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n536), .A2(new_n537), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT85), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n536), .A2(new_n533), .A3(new_n537), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n558), .A2(new_n360), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n550), .B2(new_n552), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n563), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n540), .A2(new_n554), .A3(new_n543), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(KEYINPUT88), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n561), .A2(KEYINPUT20), .A3(new_n562), .A4(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n562), .B1(new_n555), .B2(new_n560), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n543), .B1(new_n540), .B2(new_n554), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n371), .B1(new_n555), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G475), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n574), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(G234), .A2(G237), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n583), .A2(G952), .A3(new_n364), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n583), .A2(G902), .A3(G953), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT21), .B(G898), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n251), .A2(G122), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(KEYINPUT14), .ZN(new_n591));
  INV_X1    g405(.A(G122), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G116), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT14), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(KEYINPUT90), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(G116), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n590), .A2(KEYINPUT14), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n591), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G107), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n596), .A2(new_n590), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n398), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT89), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n193), .B2(G128), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n196), .A2(KEYINPUT89), .A3(G143), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n193), .A2(G128), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n205), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n205), .B1(new_n605), .B2(new_n606), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n599), .B(new_n601), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n600), .B(new_n398), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n606), .B(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n605), .ZN(new_n614));
  OAI21_X1  g428(.A(G134), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n615), .A3(new_n607), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n467), .A2(new_n379), .A3(G953), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT91), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n610), .A2(new_n619), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n371), .ZN(new_n624));
  INV_X1    g438(.A(G478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT15), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n582), .A2(new_n588), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n337), .A2(new_n389), .A3(new_n522), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  NOR2_X1   g448(.A1(new_n471), .A2(new_n388), .ZN(new_n635));
  INV_X1    g449(.A(new_n519), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n516), .B1(new_n501), .B2(new_n514), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n472), .B(new_n588), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n622), .A2(KEYINPUT33), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n619), .B1(new_n610), .B2(new_n616), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT93), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n639), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n625), .A2(G902), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT92), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n623), .B2(new_n647), .ZN(new_n648));
  AOI211_X1 g462(.A(KEYINPUT92), .B(KEYINPUT33), .C1(new_n621), .C2(new_n622), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n644), .B(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n624), .A2(new_n625), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n581), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n638), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n325), .B1(new_n316), .B2(new_n371), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n323), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n635), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  AND2_X1   g473(.A1(new_n574), .A2(new_n580), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n561), .A2(new_n573), .ZN(new_n661));
  INV_X1    g475(.A(new_n562), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n576), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n660), .A2(new_n629), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n638), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n635), .A2(new_n656), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT94), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT35), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G107), .ZN(G9));
  NOR2_X1   g483(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n363), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n386), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n383), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT95), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT95), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n383), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT96), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT96), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n382), .A2(new_n380), .ZN(new_n680));
  AOI211_X1 g494(.A(KEYINPUT95), .B(new_n672), .C1(new_n680), .C2(new_n378), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n676), .B1(new_n383), .B2(new_n673), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n522), .A2(new_n632), .A3(new_n684), .A4(new_n656), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT37), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n686), .B(KEYINPUT97), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G110), .ZN(G12));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n585), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n584), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n660), .A2(new_n629), .A3(new_n663), .A4(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n678), .B2(new_n683), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n337), .A2(new_n694), .A3(new_n522), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  INV_X1    g510(.A(new_n471), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n692), .B(KEYINPUT39), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT40), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n289), .A2(new_n306), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n283), .B1(new_n331), .B2(new_n287), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n371), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n321), .A2(new_n324), .A3(new_n701), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n518), .A2(new_n519), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT38), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n675), .A2(new_n677), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n581), .A2(new_n629), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n708), .A2(new_n709), .A3(new_n473), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n700), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NAND3_X1  g527(.A1(new_n581), .A2(new_n652), .A3(new_n692), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n678), .B2(new_n683), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n337), .A2(new_n522), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n461), .A2(new_n468), .ZN(new_n719));
  INV_X1    g533(.A(G469), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n458), .A2(new_n371), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT99), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n458), .A2(KEYINPUT99), .A3(new_n371), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(new_n654), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n337), .A3(new_n389), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT100), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(KEYINPUT100), .A3(new_n337), .A4(new_n389), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT41), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G113), .ZN(G15));
  NAND4_X1  g547(.A1(new_n337), .A2(new_n389), .A3(new_n665), .A4(new_n725), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  NAND2_X1  g549(.A1(new_n721), .A2(new_n722), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(G469), .A3(new_n724), .ZN(new_n737));
  INV_X1    g551(.A(new_n719), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n520), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n337), .A3(new_n632), .A4(new_n684), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(new_n725), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n520), .A2(new_n629), .A3(new_n581), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n587), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n332), .A2(new_n283), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n307), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT101), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n308), .A2(new_n309), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT101), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n307), .A2(new_n750), .A3(new_n746), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n655), .B1(new_n752), .B2(new_n317), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT102), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n389), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n753), .B2(new_n389), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n745), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  AND3_X1   g573(.A1(new_n581), .A2(new_n652), .A3(new_n692), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n520), .A2(new_n737), .A3(new_n760), .A4(new_n738), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n753), .A3(new_n709), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  NAND2_X1  g577(.A1(new_n466), .A2(new_n468), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n518), .A2(new_n472), .A3(new_n519), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n337), .A2(new_n389), .A3(new_n766), .A4(new_n760), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n318), .A2(new_n320), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n768), .B(new_n388), .C1(new_n769), .C2(new_n336), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n764), .A2(new_n714), .A3(new_n765), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(G131), .Z(G33));
  INV_X1    g587(.A(new_n693), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n337), .A2(new_n389), .A3(new_n774), .A4(new_n766), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(new_n652), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n777), .A2(new_n581), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n581), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT103), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n783), .B(new_n709), .C1(new_n323), .C2(new_n655), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n433), .A2(new_n418), .A3(new_n436), .A4(new_n444), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n419), .A2(new_n425), .A3(new_n432), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n230), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n436), .B1(new_n789), .B2(new_n433), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT45), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n462), .A2(new_n463), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n793), .A3(G469), .ZN(new_n794));
  NAND2_X1  g608(.A1(G469), .A2(G902), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT46), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n461), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n468), .A3(new_n698), .ZN(new_n801));
  INV_X1    g615(.A(new_n765), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n786), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT104), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n207), .ZN(G39));
  NOR4_X1   g620(.A1(new_n337), .A2(new_n389), .A3(new_n714), .A4(new_n765), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT106), .Z(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT105), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n800), .B2(new_n468), .ZN(new_n811));
  INV_X1    g625(.A(new_n468), .ZN(new_n812));
  AOI211_X1 g626(.A(KEYINPUT105), .B(new_n812), .C1(new_n798), .C2(new_n799), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n809), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n799), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n815), .A2(new_n796), .A3(new_n797), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT105), .B1(new_n816), .B2(new_n812), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n800), .A2(new_n810), .A3(new_n468), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n808), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G140), .ZN(G42));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NOR2_X1   g637(.A1(G952), .A2(G953), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT116), .Z(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n725), .A2(new_n584), .A3(new_n802), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n706), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n389), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n582), .A2(new_n777), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n783), .ZN(new_n832));
  INV_X1    g646(.A(new_n655), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n307), .A2(new_n750), .A3(new_n746), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n750), .B1(new_n307), .B2(new_n746), .ZN(new_n835));
  INV_X1    g649(.A(new_n749), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n833), .B(new_n709), .C1(new_n837), .C2(new_n322), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n830), .A2(new_n831), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n783), .A2(new_n584), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n753), .A2(new_n389), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT102), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n765), .B(new_n840), .C1(new_n842), .C2(new_n755), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n797), .B1(new_n723), .B2(new_n724), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n469), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n814), .A2(new_n819), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n839), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n725), .A2(new_n848), .A3(new_n473), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n708), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n725), .B2(new_n473), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n840), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n852), .B(new_n853), .C1(new_n756), .C2(new_n757), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT50), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n855), .B1(new_n854), .B2(KEYINPUT112), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n847), .B(KEYINPUT51), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(KEYINPUT112), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT50), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT51), .A4(new_n847), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n769), .A2(new_n336), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n389), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n832), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT48), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n830), .A2(new_n653), .ZN(new_n873));
  INV_X1    g687(.A(G952), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(G953), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n840), .B1(new_n842), .B2(new_n755), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n876), .A2(KEYINPUT114), .A3(new_n740), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT114), .B1(new_n876), .B2(new_n740), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n872), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n866), .A2(new_n867), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n867), .B1(new_n866), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n383), .A2(new_n673), .A3(new_n692), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n520), .A2(new_n886), .A3(new_n629), .A4(new_n581), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n764), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n706), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n762), .A2(new_n695), .A3(new_n716), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n741), .A2(new_n734), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n731), .A2(new_n758), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n582), .A2(new_n630), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n777), .A2(new_n581), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n638), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n635), .A3(new_n899), .A4(new_n656), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n633), .A2(new_n685), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT107), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n633), .A2(KEYINPUT107), .A3(new_n900), .A4(new_n685), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n753), .A2(new_n771), .A3(new_n709), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n660), .A2(new_n630), .A3(new_n663), .A4(new_n692), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n765), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n337), .A2(new_n697), .A3(new_n684), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n775), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n772), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n892), .A2(new_n895), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n893), .B1(new_n729), .B2(new_n730), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n905), .A2(new_n916), .A3(new_n911), .A4(new_n758), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n725), .A2(new_n520), .A3(new_n760), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n695), .B1(new_n838), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n716), .A2(new_n889), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n891), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n891), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n695), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT108), .B1(new_n762), .B2(new_n695), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT109), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n890), .A2(new_n927), .A3(new_n891), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n922), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT110), .A4(new_n928), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n917), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n915), .B1(new_n933), .B2(KEYINPUT53), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n917), .A2(new_n913), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT108), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n838), .A2(new_n918), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n337), .A2(new_n522), .A3(new_n694), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n695), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI22_X1  g755(.A1(new_n941), .A2(new_n923), .B1(new_n921), .B2(KEYINPUT109), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT110), .B1(new_n942), .B2(new_n928), .ZN(new_n943));
  AND4_X1   g757(.A1(KEYINPUT110), .A2(new_n922), .A3(new_n926), .A4(new_n928), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT54), .B1(new_n912), .B2(new_n913), .ZN(new_n946));
  AOI22_X1  g760(.A1(new_n934), .A2(KEYINPUT54), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n826), .B1(new_n885), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n388), .A2(new_n469), .A3(new_n473), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n829), .A2(new_n708), .A3(new_n780), .A4(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n844), .B(KEYINPUT49), .Z(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n823), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n866), .A2(new_n882), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT115), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n866), .A2(new_n867), .A3(new_n882), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n945), .A2(new_n946), .ZN(new_n958));
  INV_X1    g772(.A(new_n917), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n943), .B2(new_n944), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n914), .B1(new_n960), .B2(new_n913), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT54), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n825), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n952), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(KEYINPUT117), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n953), .A2(new_n966), .ZN(G75));
  XNOR2_X1  g781(.A(new_n890), .B(KEYINPUT52), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n913), .B1(new_n917), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n371), .B1(new_n945), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(G210), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT56), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n499), .A2(new_n500), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(new_n485), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT55), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n364), .A2(G952), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(G51));
  INV_X1    g793(.A(KEYINPUT118), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n905), .A4(new_n911), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n931), .B2(new_n932), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n969), .A2(new_n962), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n945), .A2(KEYINPUT118), .A3(new_n946), .ZN(new_n985));
  INV_X1    g799(.A(new_n969), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT54), .B1(new_n982), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n795), .B(KEYINPUT57), .Z(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n458), .ZN(new_n991));
  INV_X1    g805(.A(new_n794), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n970), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n978), .B1(new_n991), .B2(new_n993), .ZN(G54));
  INV_X1    g808(.A(KEYINPUT119), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n970), .A2(KEYINPUT58), .A3(G475), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n661), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n978), .B1(new_n996), .B2(new_n661), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n996), .A2(new_n995), .A3(new_n661), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(G60));
  INV_X1    g815(.A(new_n648), .ZN(new_n1002));
  INV_X1    g816(.A(new_n649), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n640), .A2(new_n643), .ZN(new_n1004));
  AOI22_X1  g818(.A1(new_n1002), .A2(new_n1003), .B1(new_n1004), .B2(new_n639), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G478), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT59), .Z(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT120), .B1(new_n988), .B2(new_n1010), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n988), .A2(KEYINPUT120), .A3(new_n1010), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1005), .B1(new_n963), .B2(new_n1008), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT121), .ZN(new_n1014));
  OAI22_X1  g828(.A1(new_n1011), .A2(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n978), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1005), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n947), .B2(new_n1007), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1018), .B2(KEYINPUT121), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1015), .A2(new_n1019), .ZN(G63));
  NAND2_X1  g834(.A1(new_n945), .A2(new_n969), .ZN(new_n1021));
  XNOR2_X1  g835(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n379), .A2(new_n371), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n385), .ZN(new_n1026));
  NOR2_X1   g840(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n978), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n671), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1026), .B(new_n1028), .C1(new_n1029), .C2(new_n1025), .ZN(new_n1030));
  NAND2_X1  g844(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1030), .B(new_n1031), .ZN(G66));
  NOR3_X1   g846(.A1(new_n586), .A2(new_n480), .A3(new_n364), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n895), .A2(new_n905), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(new_n364), .ZN(new_n1036));
  INV_X1    g850(.A(G898), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n973), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1036), .B(new_n1038), .Z(G69));
  OAI21_X1  g853(.A(new_n293), .B1(new_n262), .B2(new_n265), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n557), .B(KEYINPUT124), .Z(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G900), .A2(G953), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n869), .A2(new_n744), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n801), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1045), .B(KEYINPUT125), .ZN(new_n1046));
  INV_X1    g860(.A(new_n775), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n804), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n772), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n941), .A2(new_n716), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n1048), .A2(new_n1049), .A3(new_n821), .A4(new_n1050), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n1042), .B(new_n1043), .C1(new_n1051), .C2(G953), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1050), .A2(new_n712), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1055));
  INV_X1    g869(.A(new_n898), .ZN(new_n1056));
  NOR3_X1   g870(.A1(new_n1056), .A2(new_n699), .A3(new_n765), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1057), .A2(new_n337), .A3(new_n389), .ZN(new_n1058));
  AOI211_X1 g872(.A(new_n1058), .B(new_n804), .C1(new_n820), .C2(new_n808), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1054), .A2(new_n1055), .A3(new_n1059), .ZN(new_n1060));
  AND2_X1   g874(.A1(new_n1060), .A2(new_n364), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1052), .B1(new_n1061), .B2(new_n1042), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n364), .B1(G227), .B2(G900), .ZN(new_n1063));
  XNOR2_X1  g877(.A(new_n1062), .B(new_n1063), .ZN(G72));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n1060), .B2(new_n1034), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n328), .A2(new_n303), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g883(.A(KEYINPUT126), .ZN(new_n1070));
  XNOR2_X1  g884(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  OAI211_X1 g885(.A(new_n289), .B(new_n306), .C1(new_n283), .C2(new_n328), .ZN(new_n1072));
  NAND3_X1  g886(.A1(new_n934), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1066), .B1(new_n1051), .B2(new_n1034), .ZN(new_n1074));
  XNOR2_X1  g888(.A(new_n1074), .B(KEYINPUT127), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n328), .A2(new_n303), .ZN(new_n1076));
  OAI211_X1 g890(.A(new_n1016), .B(new_n1073), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n1071), .A2(new_n1077), .ZN(G57));
endmodule


