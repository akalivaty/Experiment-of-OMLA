//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(new_n203), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NOR2_X1   g0017(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n218));
  AND2_X1   g0018(.A1(G77), .A2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n219), .B(new_n223), .C1(G116), .C2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n218), .B1(new_n229), .B2(new_n214), .ZN(new_n230));
  NAND2_X1  g0030(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n213), .B(new_n217), .C1(new_n232), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n228), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n225), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n227), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n225), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n212), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(new_n253), .B2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT8), .A2(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT8), .A2(G58), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT69), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n211), .A2(G33), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT70), .B(new_n265), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n201), .ZN(new_n275));
  OAI21_X1  g0075(.A(G20), .B1(new_n275), .B2(new_n209), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n269), .B2(new_n271), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n264), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  AND3_X1   g0080(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n258), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT71), .B1(new_n280), .B2(new_n258), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n256), .B(new_n260), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n289), .B2(G226), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G222), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G223), .A2(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n287), .C1(G77), .C2(new_n291), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G179), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n283), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(G200), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n290), .A2(G190), .A3(new_n296), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT9), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n303), .B(new_n304), .C1(new_n283), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n283), .A2(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n311), .B2(new_n306), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n288), .A2(new_n284), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n288), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G238), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n228), .A2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G226), .B2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n319), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n286), .B1(new_n327), .B2(new_n287), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n318), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT14), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(G179), .A3(new_n332), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n337), .A3(G169), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  OAI22_X1  g0139(.A1(new_n262), .A2(new_n225), .B1(new_n211), .B2(G68), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n273), .A2(new_n202), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n258), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT74), .B(KEYINPUT11), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n254), .A2(KEYINPUT12), .A3(G68), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT12), .B1(new_n254), .B2(G68), .ZN(new_n346));
  AOI22_X1  g0146(.A1(G68), .A2(new_n259), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n258), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT7), .B1(new_n326), .B2(new_n211), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  AOI211_X1 g0152(.A(new_n352), .B(G20), .C1(new_n323), .C2(new_n325), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G68), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n227), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n203), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n261), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT16), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n354), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n272), .A2(new_n254), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n272), .A2(new_n259), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n363), .A2(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n226), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n323), .A2(new_n368), .A3(new_n325), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n287), .ZN(new_n373));
  INV_X1    g0173(.A(new_n286), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n288), .A2(G232), .A3(new_n284), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G200), .ZN(new_n377));
  INV_X1    g0177(.A(G190), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n367), .A2(KEYINPUT17), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n352), .B1(new_n291), .B2(G20), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n324), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n383));
  OAI211_X1 g0183(.A(KEYINPUT7), .B(new_n211), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n355), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n362), .B1(new_n385), .B2(new_n359), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n364), .A2(new_n386), .A3(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n366), .A2(new_n365), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n379), .A3(new_n377), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n380), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n388), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n376), .A2(G169), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n373), .A2(G179), .A3(new_n374), .A4(new_n375), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT18), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  AOI221_X4 g0198(.A(new_n398), .B1(new_n394), .B2(new_n395), .C1(new_n387), .C2(new_n388), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(KEYINPUT75), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n393), .A2(KEYINPUT18), .A3(new_n396), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n392), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n333), .A2(G200), .ZN(new_n405));
  INV_X1    g0205(.A(new_n348), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(new_n406), .C1(new_n378), .C2(new_n333), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n286), .B1(new_n289), .B2(G244), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G238), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n291), .B(new_n409), .C1(new_n228), .C2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n287), .C1(G107), .C2(new_n291), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n412), .A2(G169), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n254), .A2(G77), .ZN(new_n414));
  INV_X1    g0214(.A(new_n268), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n261), .B1(G20), .B2(G77), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT15), .B(G87), .Z(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(new_n273), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n414), .B1(new_n419), .B2(new_n258), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n259), .A2(G77), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n412), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AND4_X1   g0225(.A1(new_n349), .A2(new_n404), .A3(new_n407), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n412), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT72), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n412), .A2(G190), .ZN(new_n430));
  INV_X1    g0230(.A(new_n421), .ZN(new_n431));
  AOI211_X1 g0231(.A(new_n414), .B(new_n431), .C1(new_n419), .C2(new_n258), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n432), .B(new_n433), .C1(new_n427), .C2(new_n412), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n313), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G303), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n326), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G264), .A2(G1698), .ZN(new_n439));
  INV_X1    g0239(.A(G257), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(new_n287), .C1(new_n326), .C2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n253), .A2(G45), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(new_n285), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n288), .A3(G270), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n442), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT78), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n442), .A2(new_n447), .A3(new_n451), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G190), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n253), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n350), .A2(new_n455), .A3(new_n254), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n254), .A2(G116), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT79), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n211), .C1(G33), .C2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n258), .C1(new_n211), .C2(G116), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n458), .B(new_n460), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n454), .B(new_n469), .C1(new_n427), .C2(new_n453), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n468), .A2(new_n450), .A3(G169), .A4(new_n452), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT21), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n449), .A2(new_n423), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n468), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n470), .A2(new_n473), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n471), .B(KEYINPUT21), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n476), .A4(new_n470), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n291), .A2(G244), .A3(new_n292), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT77), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(KEYINPUT77), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n291), .A2(G250), .A3(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n461), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n287), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n446), .A2(new_n288), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(G257), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n447), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n462), .A2(new_n496), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(new_n206), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(KEYINPUT6), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(G20), .B1(G77), .B2(new_n261), .ZN(new_n501));
  OAI21_X1  g0301(.A(G107), .B1(new_n351), .B2(new_n353), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n350), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n456), .A2(new_n462), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n255), .A2(new_n462), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT76), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n495), .B(new_n507), .C1(new_n378), .C2(new_n494), .ZN(new_n508));
  INV_X1    g0308(.A(new_n447), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n509), .B(new_n492), .C1(new_n489), .C2(new_n287), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n423), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n494), .A2(new_n299), .ZN(new_n512));
  INV_X1    g0312(.A(new_n507), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n292), .A2(G244), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n291), .B(new_n515), .C1(G238), .C2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G116), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n288), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n443), .A2(G250), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n287), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n443), .A2(new_n285), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT19), .B1(new_n207), .B2(G87), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n211), .B2(new_n319), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n291), .A2(new_n211), .A3(G68), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n319), .A2(G20), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(KEYINPUT19), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n258), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n418), .A2(new_n255), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n457), .A2(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n520), .A2(new_n521), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n516), .A2(new_n517), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n288), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n523), .A2(new_n531), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n529), .B(new_n530), .C1(new_n456), .C2(new_n418), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n522), .A2(new_n423), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(new_n299), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n508), .A2(new_n514), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(G250), .A2(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n440), .A2(G1698), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n323), .A2(new_n544), .A3(new_n325), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT81), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(KEYINPUT81), .A3(new_n547), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(new_n287), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n491), .A2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n447), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n427), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n378), .A3(new_n447), .A4(new_n553), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n457), .A2(G107), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n254), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n323), .A2(new_n325), .A3(new_n211), .A4(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n291), .A2(new_n563), .A3(new_n211), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n211), .A2(G107), .ZN(new_n566));
  XNOR2_X1  g0366(.A(new_n566), .B(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n565), .A2(KEYINPUT24), .A3(new_n567), .A4(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n258), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n557), .A2(new_n558), .A3(new_n560), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n558), .A3(new_n560), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n554), .A2(G179), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n554), .A2(new_n299), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT82), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n574), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n482), .A2(new_n543), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n436), .A2(new_n584), .ZN(G372));
  NOR2_X1   g0385(.A1(new_n399), .A2(new_n397), .ZN(new_n586));
  INV_X1    g0386(.A(new_n425), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n407), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n349), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n389), .B(KEYINPUT17), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n591), .A2(new_n592), .B1(new_n312), .B2(new_n310), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n302), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n574), .A2(new_n508), .A3(new_n514), .A4(new_n542), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT83), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n480), .A2(new_n476), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n541), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n511), .A2(new_n512), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT26), .A3(new_n513), .A4(new_n542), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n537), .A2(new_n541), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n514), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n595), .B1(new_n436), .B2(new_n609), .ZN(G369));
  INV_X1    g0410(.A(G13), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n253), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(G213), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G343), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n575), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n574), .A2(new_n578), .A3(new_n581), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n581), .B1(new_n574), .B2(new_n578), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n625));
  INV_X1    g0425(.A(new_n618), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(new_n625), .C1(new_n578), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n482), .B1(new_n469), .B2(new_n626), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n469), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n599), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G330), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n598), .A2(new_n626), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n625), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n599), .A2(new_n626), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(G399));
  INV_X1    g0442(.A(new_n215), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G1), .ZN(new_n646));
  INV_X1    g0446(.A(G87), .ZN(new_n647));
  INV_X1    g0447(.A(G116), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n462), .A3(new_n496), .A4(new_n648), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n646), .A2(new_n649), .B1(new_n210), .B2(new_n645), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  AOI211_X1 g0451(.A(KEYINPUT29), .B(new_n618), .C1(new_n600), .C2(new_n607), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n607), .A2(KEYINPUT86), .ZN(new_n653));
  OR3_X1    g0453(.A1(new_n599), .A2(KEYINPUT87), .A3(new_n597), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT87), .B1(new_n599), .B2(new_n597), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n596), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n607), .A2(KEYINPUT86), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n626), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n659), .B2(KEYINPUT29), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n482), .A2(new_n543), .A3(new_n583), .A4(new_n626), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT30), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n490), .A2(new_n447), .A3(new_n493), .A4(new_n522), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n475), .A2(new_n553), .A3(new_n552), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n552), .A2(new_n553), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n666), .A2(new_n423), .A3(new_n449), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n522), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n494), .A2(new_n423), .A3(new_n554), .A4(new_n535), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n665), .B(new_n668), .C1(new_n669), .C2(new_n453), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n618), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT31), .B1(new_n670), .B2(new_n618), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n661), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n651), .B1(new_n676), .B2(G1), .ZN(G364));
  AOI21_X1  g0477(.A(new_n646), .B1(G45), .B2(new_n612), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n632), .ZN(new_n680));
  NOR2_X1   g0480(.A1(G13), .A2(G33), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n211), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT93), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n212), .B1(G20), .B2(new_n299), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n378), .A2(G179), .A3(G200), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n211), .ZN(new_n688));
  INV_X1    g0488(.A(G294), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n211), .A2(G190), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(new_n423), .A3(new_n427), .ZN(new_n691));
  INV_X1    g0491(.A(G329), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n688), .A2(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n423), .A2(G200), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT90), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n211), .A2(new_n378), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n291), .B1(new_n698), .B2(G303), .ZN(new_n699));
  INV_X1    g0499(.A(G283), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n690), .ZN(new_n701));
  INV_X1    g0501(.A(G311), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n423), .A2(G200), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n690), .ZN(new_n704));
  OAI221_X1 g0504(.A(new_n699), .B1(new_n700), .B2(new_n701), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n423), .A2(new_n427), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n690), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g0508(.A(KEYINPUT33), .B(G317), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n693), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G322), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n696), .A2(new_n703), .ZN(new_n712));
  INV_X1    g0512(.A(G326), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n696), .A2(new_n706), .ZN(new_n714));
  OAI221_X1 g0514(.A(new_n710), .B1(new_n711), .B2(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n697), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n326), .B1(new_n716), .B2(G87), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(KEYINPUT91), .ZN(new_n718));
  INV_X1    g0518(.A(new_n712), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(G58), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n701), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G107), .ZN(new_n722));
  INV_X1    g0522(.A(new_n714), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G50), .ZN(new_n724));
  INV_X1    g0524(.A(new_n691), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G159), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT89), .B(KEYINPUT32), .Z(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n726), .A2(new_n727), .B1(G68), .B2(new_n708), .ZN(new_n729));
  INV_X1    g0529(.A(new_n688), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G97), .ZN(new_n731));
  INV_X1    g0531(.A(new_n704), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G77), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n728), .A2(new_n729), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(KEYINPUT91), .B2(new_n717), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n720), .A2(new_n722), .A3(new_n724), .A4(new_n735), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n715), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n682), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n685), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n251), .A2(G45), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n326), .A2(new_n215), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT88), .Z(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n210), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n741), .A2(new_n744), .B1(G116), .B2(new_n215), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n643), .A2(new_n326), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(G355), .B2(new_n746), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n684), .B1(new_n686), .B2(new_n737), .C1(new_n740), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n632), .A2(G330), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n633), .A2(new_n679), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(G396));
  AOI21_X1  g0551(.A(new_n618), .B1(new_n600), .B2(new_n607), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n435), .B1(new_n432), .B2(new_n626), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n425), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n587), .A2(new_n626), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n752), .B(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n679), .B1(new_n758), .B2(new_n675), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT96), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n758), .A2(new_n675), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n714), .A2(new_n437), .B1(new_n704), .B2(new_n648), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(G283), .B2(new_n708), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  AOI21_X1  g0565(.A(new_n291), .B1(new_n698), .B2(G107), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT95), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n730), .A2(G97), .B1(new_n725), .B2(G311), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n647), .C2(new_n701), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n765), .B(new_n769), .C1(G294), .C2(new_n719), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G143), .A2(new_n719), .B1(new_n708), .B2(G150), .ZN(new_n771));
  INV_X1    g0571(.A(G137), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n771), .B1(new_n772), .B2(new_n714), .C1(new_n773), .C2(new_n704), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT34), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n774), .A2(new_n775), .B1(G58), .B2(new_n730), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n721), .A2(G68), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n326), .B1(new_n698), .B2(G50), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n776), .B(new_n780), .C1(G132), .C2(new_n725), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n685), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n685), .A2(new_n681), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n202), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n756), .A2(new_n681), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n782), .A2(new_n678), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n762), .A2(new_n786), .ZN(G384));
  AND2_X1   g0587(.A1(new_n339), .A2(new_n348), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n626), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT101), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT39), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT38), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n393), .A2(new_n396), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n398), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n393), .A2(KEYINPUT75), .A3(KEYINPUT18), .A4(new_n396), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n403), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n590), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT97), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(KEYINPUT16), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n258), .B1(new_n361), .B2(new_n799), .C1(new_n798), .C2(new_n386), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n388), .ZN(new_n801));
  INV_X1    g0601(.A(new_n616), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(KEYINPUT98), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT98), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n806), .B(new_n803), .C1(new_n796), .C2(new_n590), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT37), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n801), .B1(new_n396), .B2(new_n802), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n389), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT99), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n393), .A2(new_n812), .A3(new_n396), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n393), .A2(new_n802), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n813), .A2(new_n814), .A3(new_n809), .A4(new_n389), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n812), .B1(new_n393), .B2(new_n396), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT100), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT100), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n815), .B2(new_n816), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n811), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n792), .B1(new_n808), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n811), .ZN(new_n823));
  INV_X1    g0623(.A(new_n820), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n826), .B(KEYINPUT38), .C1(new_n805), .C2(new_n807), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n791), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n814), .A2(new_n389), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n809), .B1(new_n829), .B2(new_n793), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n818), .B2(new_n820), .ZN(new_n831));
  INV_X1    g0631(.A(new_n586), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n814), .B1(new_n832), .B2(new_n590), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n792), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n827), .A2(new_n791), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT102), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n827), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n806), .B1(new_n404), .B2(new_n803), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n797), .A2(KEYINPUT98), .A3(new_n804), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT38), .B1(new_n840), .B2(new_n826), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT39), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT102), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n827), .A2(new_n834), .A3(new_n791), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n790), .B1(new_n836), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n837), .A2(new_n841), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n755), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n752), .B2(new_n754), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n349), .B(new_n407), .C1(new_n406), .C2(new_n626), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n788), .A2(new_n618), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n848), .A2(new_n855), .B1(new_n586), .B2(new_n616), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n827), .A2(new_n834), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n756), .B1(new_n851), .B2(new_n852), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(KEYINPUT40), .A3(new_n674), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n674), .A2(new_n860), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n822), .B2(new_n827), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(G330), .C1(new_n863), .C2(KEYINPUT40), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n436), .A2(new_n675), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n847), .B2(new_n862), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n674), .A3(new_n861), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n436), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n858), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n595), .B1(new_n660), .B2(new_n436), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n253), .B2(new_n612), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n648), .B1(new_n500), .B2(KEYINPUT35), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n212), .A2(new_n211), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(KEYINPUT35), .C2(new_n500), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n210), .A2(new_n202), .A3(new_n356), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n275), .A2(new_n355), .ZN(new_n881));
  OAI211_X1 g0681(.A(G1), .B(new_n611), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n875), .A2(new_n879), .A3(new_n882), .ZN(G367));
  NAND2_X1  g0683(.A1(new_n513), .A2(new_n618), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n508), .A2(new_n514), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n602), .A2(new_n513), .A3(new_n618), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n635), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT103), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT42), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n639), .B1(new_n623), .B2(new_n625), .ZN(new_n891));
  INV_X1    g0691(.A(new_n887), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n885), .A2(new_n578), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n618), .B1(new_n894), .B2(new_n514), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n889), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n639), .B(new_n887), .C1(new_n623), .C2(new_n625), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n890), .ZN(new_n898));
  INV_X1    g0698(.A(new_n895), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT103), .B(new_n899), .C1(new_n897), .C2(new_n890), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n531), .A2(new_n532), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n618), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n542), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n601), .A2(new_n902), .A3(new_n618), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT43), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n910));
  INV_X1    g0710(.A(new_n906), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n907), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n901), .A2(new_n914), .A3(new_n908), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n910), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT105), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n910), .A2(new_n913), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n888), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n253), .B1(new_n612), .B2(G45), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT45), .B1(new_n641), .B2(new_n892), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT45), .ZN(new_n925));
  NOR4_X1   g0725(.A1(new_n891), .A2(new_n925), .A3(new_n637), .A4(new_n887), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n641), .B2(new_n892), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n887), .B(new_n928), .C1(new_n891), .C2(new_n637), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n634), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n624), .B1(new_n583), .B2(new_n619), .ZN(new_n934));
  INV_X1    g0734(.A(new_n625), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n640), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n636), .A3(new_n892), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n925), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n641), .A2(KEYINPUT45), .A3(new_n892), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n940), .A2(new_n635), .A3(new_n931), .A4(new_n930), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n936), .B1(new_n627), .B2(new_n640), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(new_n633), .Z(new_n943));
  NAND4_X1  g0743(.A1(new_n933), .A2(new_n676), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n676), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n644), .B(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n923), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n917), .A2(new_n888), .A3(new_n919), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n921), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n291), .B1(new_n712), .B2(new_n263), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n721), .A2(G77), .B1(G137), .B2(new_n725), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n355), .B2(new_n688), .C1(new_n201), .C2(new_n704), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(G143), .C2(new_n723), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n227), .B2(new_n697), .C1(new_n773), .C2(new_n707), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n714), .A2(new_n702), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n725), .A2(G317), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n697), .A2(new_n648), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n957), .B1(new_n496), .B2(new_n688), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(KEYINPUT46), .A2(G116), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n698), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n701), .A2(new_n462), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n437), .B2(new_n712), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G294), .B2(new_n708), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n732), .A2(G283), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n962), .A2(new_n966), .A3(new_n326), .A4(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n955), .B1(new_n956), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n685), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n911), .A2(new_n683), .ZN(new_n972));
  INV_X1    g0772(.A(new_n743), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n739), .B1(new_n215), .B2(new_n418), .C1(new_n242), .C2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n971), .A2(new_n678), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n950), .A2(new_n975), .ZN(G387));
  OR2_X1    g0776(.A1(new_n676), .A2(new_n943), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n676), .A2(new_n943), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n644), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n326), .B1(new_n691), .B2(new_n713), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G311), .A2(new_n708), .B1(new_n719), .B2(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n437), .B2(new_n704), .C1(new_n711), .C2(new_n714), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n700), .B2(new_n688), .C1(new_n689), .C2(new_n697), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT49), .Z(new_n985));
  AOI211_X1 g0785(.A(new_n980), .B(new_n985), .C1(G116), .C2(new_n721), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n272), .A2(new_n707), .B1(new_n355), .B2(new_n704), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT108), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n714), .A2(new_n773), .B1(new_n712), .B2(new_n225), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n418), .A2(new_n688), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(G150), .C2(new_n725), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n964), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n697), .A2(new_n202), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n992), .A2(new_n326), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n685), .B1(new_n986), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n679), .B1(new_n628), .B2(new_n683), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n973), .B1(new_n238), .B2(G45), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n649), .B2(new_n746), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n415), .A2(new_n225), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n355), .A2(new_n202), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n1001), .A2(G45), .A3(new_n1002), .A4(new_n649), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n999), .A2(new_n1003), .B1(G107), .B2(new_n215), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n997), .B1(new_n739), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n943), .B2(new_n923), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n979), .A2(new_n1006), .ZN(G393));
  INV_X1    g0807(.A(KEYINPUT109), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n933), .A2(new_n1008), .A3(new_n941), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n927), .A2(new_n932), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT109), .A3(new_n635), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n978), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1009), .A2(new_n1011), .A3(new_n1014), .A4(new_n978), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1013), .A2(new_n644), .A3(new_n944), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n887), .A2(new_n738), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n714), .A2(new_n1019), .B1(new_n712), .B2(new_n702), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT52), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n291), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n722), .B1(new_n700), .B2(new_n697), .C1(new_n689), .C2(new_n704), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G116), .C2(new_n730), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n437), .B2(new_n707), .C1(new_n711), .C2(new_n691), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n688), .A2(new_n202), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n701), .A2(new_n647), .B1(new_n268), .B2(new_n704), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G68), .C2(new_n716), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n725), .A2(G143), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n708), .A2(new_n275), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n714), .A2(new_n263), .B1(new_n712), .B2(new_n773), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT51), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n326), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n686), .B1(new_n1027), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n215), .A2(new_n462), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n740), .B(new_n1040), .C1(new_n248), .C2(new_n743), .ZN(new_n1041));
  OR4_X1    g0841(.A1(new_n679), .A2(new_n1018), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n923), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1016), .A2(new_n1042), .A3(new_n1044), .ZN(G390));
  OAI21_X1  g0845(.A(new_n790), .B1(new_n850), .B2(new_n854), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n836), .A2(new_n845), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT86), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n607), .B(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n618), .B1(new_n1049), .B2(new_n656), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n849), .B1(new_n1050), .B2(new_n754), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n790), .B(new_n859), .C1(new_n1051), .C2(new_n854), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n675), .A2(new_n756), .A3(new_n854), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n1047), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1054), .B1(new_n1047), .B2(new_n1052), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n866), .B(new_n595), .C1(new_n660), .C2(new_n436), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n850), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n675), .A2(new_n756), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1060), .A2(new_n853), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1061), .B2(new_n1053), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT112), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n854), .B1(new_n1063), .B2(new_n756), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n1051), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1058), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n645), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1055), .A2(new_n1056), .A3(new_n922), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n836), .A2(new_n845), .A3(new_n681), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n707), .A2(new_n496), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1028), .B1(G116), .B2(new_n719), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n700), .B2(new_n714), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G97), .B2(new_n732), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n291), .B1(new_n698), .B2(G87), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n778), .A3(new_n1079), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1075), .B(new_n1080), .C1(G294), .C2(new_n725), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n326), .B1(new_n721), .B2(new_n275), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n708), .A2(G137), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n730), .A2(G159), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  AOI22_X1  g0885(.A1(G128), .A2(new_n723), .B1(new_n732), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT53), .B1(new_n697), .B2(new_n263), .ZN(new_n1088));
  INV_X1    g0888(.A(G132), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n712), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n725), .A2(G125), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n697), .A2(KEYINPUT53), .A3(new_n263), .ZN(new_n1092));
  NOR4_X1   g0892(.A1(new_n1087), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n685), .B1(new_n1081), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1074), .A2(new_n678), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n272), .B2(new_n783), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1073), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1072), .A2(new_n1097), .ZN(G378));
  NAND2_X1  g0898(.A1(new_n283), .A2(new_n802), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT118), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n313), .A2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(KEYINPUT118), .B(new_n302), .C1(new_n310), .C2(new_n312), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n311), .A2(new_n306), .A3(KEYINPUT10), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n301), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n313), .A2(new_n1103), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n1101), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1106), .A2(new_n1112), .A3(new_n681), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(G33), .A2(G41), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT113), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n225), .C1(G41), .C2(new_n291), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n719), .A2(G128), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n707), .A2(new_n1089), .B1(new_n704), .B2(new_n772), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT115), .Z(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G125), .C2(new_n723), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n263), .B2(new_n688), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n716), .B2(new_n1085), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT59), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1115), .ZN(new_n1124));
  INV_X1    g0924(.A(G124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n725), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1128), .C1(new_n701), .C2(new_n773), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1116), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n721), .A2(G58), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT114), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n730), .A2(G68), .B1(new_n725), .B2(G283), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n462), .B2(new_n707), .C1(new_n648), .C2(new_n714), .ZN(new_n1134));
  AOI211_X1 g0934(.A(G41), .B(new_n291), .C1(new_n732), .C2(new_n417), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n496), .B2(new_n712), .ZN(new_n1136));
  NOR4_X1   g0936(.A1(new_n1132), .A2(new_n1134), .A3(new_n993), .A4(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT58), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n685), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n679), .B1(new_n201), .B2(new_n783), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1113), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT120), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n790), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n828), .A2(new_n835), .A3(KEYINPUT102), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1106), .A2(new_n1112), .A3(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n869), .A2(new_n1150), .A3(G330), .A4(new_n861), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1106), .A2(new_n1112), .A3(new_n1149), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n864), .A2(new_n1152), .ZN(new_n1153));
  AND4_X1   g0953(.A1(new_n1148), .A2(new_n856), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1148), .A2(new_n856), .B1(new_n1153), .B2(new_n1151), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n864), .A2(new_n1152), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n864), .A2(new_n1152), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1157), .A2(new_n1158), .B1(new_n846), .B2(new_n857), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1148), .A2(new_n856), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(KEYINPUT120), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1143), .B1(new_n1162), .B2(new_n923), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1053), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1047), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1068), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1058), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1058), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT57), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n644), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1163), .B1(new_n1170), .B2(new_n1173), .ZN(G375));
  NAND3_X1  g0974(.A1(new_n1067), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1070), .A2(new_n946), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n922), .B1(new_n1067), .B2(new_n1062), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n783), .A2(new_n355), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n853), .A2(G13), .A3(G33), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1132), .B1(G128), .B2(new_n725), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n732), .A2(G150), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n730), .A2(G50), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n326), .B1(new_n698), .B2(G159), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT121), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n708), .A2(new_n1085), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n719), .A2(G137), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n723), .A2(G132), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n326), .B1(new_n648), .B2(new_n707), .C1(new_n701), .C2(new_n202), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n990), .B1(G283), .B2(new_n719), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n689), .B2(new_n714), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G97), .C2(new_n698), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n496), .B2(new_n704), .C1(new_n437), .C2(new_n691), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n686), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1179), .A2(new_n1195), .A3(new_n679), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1177), .B1(new_n1178), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1176), .A2(new_n1197), .ZN(G381));
  NOR4_X1   g0998(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1199));
  INV_X1    g0999(.A(G384), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  INV_X1    g1001(.A(G381), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(G407));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n617), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(G407), .A2(G213), .A3(new_n1204), .ZN(G409));
  OAI211_X1 g1005(.A(G378), .B(new_n1163), .C1(new_n1170), .C2(new_n1173), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1159), .A2(KEYINPUT120), .A3(new_n1160), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT120), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1169), .B(new_n946), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n923), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1142), .A3(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1073), .B(new_n1096), .C1(new_n1069), .C2(new_n1071), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n617), .A2(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n645), .B1(new_n1175), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n1070), .C1(new_n1216), .C2(new_n1175), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1197), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G384), .A2(new_n1197), .A3(new_n1218), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1214), .A2(new_n1215), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1224), .B(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n617), .A2(G213), .A3(G2897), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1222), .B(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT61), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1016), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n917), .A2(new_n888), .A3(new_n919), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1233), .A2(new_n920), .A3(new_n947), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n975), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1232), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n950), .A2(new_n975), .A3(G390), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(KEYINPUT123), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(G393), .B(G396), .Z(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G387), .A2(new_n1240), .A3(new_n1232), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1236), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1239), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G387), .A2(KEYINPUT124), .A3(new_n1232), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n950), .A2(new_n1249), .A3(G390), .A4(new_n975), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1242), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1231), .A2(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1206), .A2(new_n1213), .B1(G213), .B2(new_n617), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1223), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1252), .A2(new_n1230), .A3(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(KEYINPUT122), .B(KEYINPUT63), .C1(new_n1255), .C2(new_n1223), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT122), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT63), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1224), .B2(new_n1260), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1257), .A2(KEYINPUT126), .A3(new_n1258), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT126), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1252), .A2(new_n1230), .A3(new_n1256), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1254), .B1(new_n1262), .B2(new_n1266), .ZN(G405));
  XNOR2_X1  g1067(.A(G375), .B(G378), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1222), .A2(KEYINPUT127), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1222), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(new_n1252), .ZN(G402));
endmodule


