

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n722, n723, n724, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757;

  INV_X1 U376 ( .A(n726), .ZN(n357) );
  INV_X1 U377 ( .A(n726), .ZN(n360) );
  BUF_X1 U378 ( .A(n641), .Z(n356) );
  OR2_X1 U379 ( .A1(n397), .A2(n625), .ZN(n370) );
  XNOR2_X1 U380 ( .A(n572), .B(KEYINPUT109), .ZN(n752) );
  XNOR2_X1 U381 ( .A(G143), .B(n355), .ZN(n538) );
  BUF_X1 U382 ( .A(G113), .Z(n355) );
  INV_X1 U383 ( .A(G146), .ZN(n442) );
  INV_X2 U384 ( .A(G143), .ZN(n478) );
  XNOR2_X1 U385 ( .A(n420), .B(G116), .ZN(n419) );
  INV_X1 U386 ( .A(G113), .ZN(n420) );
  XNOR2_X1 U387 ( .A(n520), .B(n519), .ZN(n393) );
  NOR2_X2 U388 ( .A1(n630), .A2(n659), .ZN(n663) );
  AND2_X1 U389 ( .A1(n358), .A2(n357), .ZN(G63) );
  XNOR2_X1 U390 ( .A(n719), .B(n359), .ZN(n358) );
  INV_X1 U391 ( .A(n720), .ZN(n359) );
  XOR2_X2 U392 ( .A(G146), .B(G125), .Z(n517) );
  XNOR2_X2 U393 ( .A(n460), .B(KEYINPUT35), .ZN(n751) );
  AND2_X1 U394 ( .A1(n361), .A2(n360), .ZN(G66) );
  XNOR2_X1 U395 ( .A(n723), .B(n362), .ZN(n361) );
  INV_X1 U396 ( .A(n724), .ZN(n362) );
  XOR2_X1 U397 ( .A(G104), .B(G107), .Z(n487) );
  NOR2_X1 U398 ( .A1(n567), .A2(n568), .ZN(n686) );
  INV_X1 U399 ( .A(G953), .ZN(n743) );
  NOR2_X1 U400 ( .A1(n567), .A2(n550), .ZN(n650) );
  XNOR2_X2 U401 ( .A(n448), .B(n447), .ZN(n753) );
  XNOR2_X2 U402 ( .A(n487), .B(n486), .ZN(n396) );
  XNOR2_X2 U403 ( .A(G137), .B(n522), .ZN(n480) );
  XNOR2_X2 U404 ( .A(n521), .B(n479), .ZN(n384) );
  XNOR2_X2 U405 ( .A(n478), .B(G128), .ZN(n521) );
  XNOR2_X1 U406 ( .A(n672), .B(n385), .ZN(n619) );
  XNOR2_X1 U407 ( .A(n437), .B(n436), .ZN(n550) );
  NOR2_X1 U408 ( .A1(G902), .A2(n709), .ZN(n495) );
  INV_X1 U409 ( .A(G122), .ZN(n425) );
  BUF_X1 U410 ( .A(n713), .Z(n722) );
  AND2_X1 U411 ( .A1(n581), .A2(n441), .ZN(n440) );
  NOR2_X1 U412 ( .A1(n617), .A2(n611), .ZN(n645) );
  XNOR2_X1 U413 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U414 ( .A(n715), .B(n714), .ZN(n716) );
  OR2_X1 U415 ( .A1(n632), .A2(G902), .ZN(n380) );
  XNOR2_X1 U416 ( .A(n740), .B(n492), .ZN(n709) );
  XNOR2_X1 U417 ( .A(n411), .B(n518), .ZN(n410) );
  XNOR2_X1 U418 ( .A(n443), .B(G101), .ZN(n516) );
  XNOR2_X1 U419 ( .A(n425), .B(KEYINPUT16), .ZN(n394) );
  XNOR2_X1 U420 ( .A(n517), .B(n432), .ZN(n741) );
  INV_X1 U421 ( .A(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U422 ( .A(G131), .B(G140), .ZN(n542) );
  AND2_X2 U423 ( .A1(n450), .A2(n449), .ZN(n713) );
  XNOR2_X1 U424 ( .A(n389), .B(n388), .ZN(n377) );
  XNOR2_X2 U425 ( .A(n383), .B(KEYINPUT19), .ZN(n598) );
  XNOR2_X2 U426 ( .A(n601), .B(KEYINPUT33), .ZN(n682) );
  NOR2_X2 U427 ( .A1(n619), .A2(n623), .ZN(n601) );
  XNOR2_X2 U428 ( .A(n599), .B(n372), .ZN(n400) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT15), .ZN(n629) );
  XNOR2_X1 U430 ( .A(n493), .B(G469), .ZN(n494) );
  INV_X1 U431 ( .A(KEYINPUT85), .ZN(n452) );
  XNOR2_X1 U432 ( .A(n587), .B(n403), .ZN(n683) );
  INV_X1 U433 ( .A(KEYINPUT38), .ZN(n403) );
  NOR2_X1 U434 ( .A1(n684), .A2(n455), .ZN(n454) );
  XNOR2_X1 U435 ( .A(n541), .B(n467), .ZN(n466) );
  INV_X1 U436 ( .A(KEYINPUT95), .ZN(n467) );
  INV_X1 U437 ( .A(n542), .ZN(n541) );
  XNOR2_X1 U438 ( .A(n610), .B(n609), .ZN(n408) );
  NAND2_X1 U439 ( .A1(n445), .A2(n515), .ZN(n570) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n515) );
  AND2_X1 U441 ( .A1(n620), .A2(n446), .ZN(n445) );
  INV_X1 U442 ( .A(KEYINPUT30), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n381), .B(KEYINPUT81), .ZN(n581) );
  NAND2_X1 U444 ( .A1(n382), .A2(n573), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n752), .B(KEYINPUT83), .ZN(n382) );
  AND2_X1 U446 ( .A1(n754), .A2(n367), .ZN(n441) );
  XNOR2_X1 U447 ( .A(n563), .B(n417), .ZN(n416) );
  OR2_X1 U448 ( .A1(G237), .A2(G902), .ZN(n526) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n439) );
  NAND2_X1 U450 ( .A1(n390), .A2(n413), .ZN(n389) );
  AND2_X1 U451 ( .A1(n753), .A2(n414), .ZN(n413) );
  NOR2_X1 U452 ( .A1(n641), .A2(n653), .ZN(n397) );
  XOR2_X1 U453 ( .A(KEYINPUT106), .B(KEYINPUT9), .Z(n528) );
  XNOR2_X1 U454 ( .A(G116), .B(KEYINPUT105), .ZN(n527) );
  XNOR2_X1 U455 ( .A(n421), .B(KEYINPUT75), .ZN(n540) );
  NAND2_X1 U456 ( .A1(n743), .A2(n422), .ZN(n421) );
  INV_X1 U457 ( .A(G237), .ZN(n422) );
  NAND2_X1 U458 ( .A1(n650), .A2(n434), .ZN(n582) );
  INV_X1 U459 ( .A(n575), .ZN(n435) );
  NAND2_X1 U460 ( .A1(n418), .A2(n375), .ZN(n450) );
  NAND2_X1 U461 ( .A1(n404), .A2(n458), .ZN(n587) );
  AND2_X1 U462 ( .A1(n622), .A2(n575), .ZN(n557) );
  INV_X1 U463 ( .A(n550), .ZN(n568) );
  XNOR2_X1 U464 ( .A(n489), .B(n428), .ZN(n492) );
  XNOR2_X1 U465 ( .A(n490), .B(n488), .ZN(n428) );
  NOR2_X1 U466 ( .A1(G952), .A2(n743), .ZN(n726) );
  NAND2_X1 U467 ( .A1(n364), .A2(n465), .ZN(n464) );
  NOR2_X1 U468 ( .A1(n700), .A2(n373), .ZN(n465) );
  INV_X1 U469 ( .A(KEYINPUT82), .ZN(n417) );
  NOR2_X2 U470 ( .A1(n751), .A2(n645), .ZN(n390) );
  NAND2_X1 U471 ( .A1(n412), .A2(G224), .ZN(n411) );
  INV_X1 U472 ( .A(G953), .ZN(n412) );
  NAND2_X1 U473 ( .A1(G234), .A2(G237), .ZN(n469) );
  INV_X1 U474 ( .A(n457), .ZN(n455) );
  XNOR2_X1 U475 ( .A(G131), .B(KEYINPUT5), .ZN(n481) );
  XOR2_X1 U476 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n482) );
  XNOR2_X1 U477 ( .A(KEYINPUT3), .B(G119), .ZN(n475) );
  INV_X1 U478 ( .A(KEYINPUT70), .ZN(n388) );
  INV_X1 U479 ( .A(KEYINPUT65), .ZN(n443) );
  INV_X1 U480 ( .A(n556), .ZN(n446) );
  OR2_X1 U481 ( .A1(n672), .A2(n684), .ZN(n379) );
  NAND2_X1 U482 ( .A1(n363), .A2(n525), .ZN(n457) );
  OR2_X1 U483 ( .A1(n525), .A2(n363), .ZN(n456) );
  NOR2_X1 U484 ( .A1(n556), .A2(n555), .ZN(n575) );
  AND2_X1 U485 ( .A1(n657), .A2(n591), .ZN(n592) );
  XNOR2_X1 U486 ( .A(G137), .B(G128), .ZN(n501) );
  INV_X1 U487 ( .A(KEYINPUT10), .ZN(n432) );
  XNOR2_X1 U488 ( .A(G140), .B(KEYINPUT24), .ZN(n496) );
  XOR2_X1 U489 ( .A(KEYINPUT97), .B(KEYINPUT23), .Z(n497) );
  XNOR2_X1 U490 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n499) );
  INV_X1 U491 ( .A(G134), .ZN(n479) );
  XNOR2_X1 U492 ( .A(G122), .B(G107), .ZN(n530) );
  XNOR2_X1 U493 ( .A(n423), .B(n544), .ZN(n546) );
  XNOR2_X1 U494 ( .A(n543), .B(n424), .ZN(n423) );
  INV_X1 U495 ( .A(KEYINPUT11), .ZN(n424) );
  XOR2_X1 U496 ( .A(G104), .B(G122), .Z(n539) );
  XNOR2_X1 U497 ( .A(KEYINPUT90), .B(G110), .ZN(n486) );
  INV_X1 U498 ( .A(KEYINPUT96), .ZN(n395) );
  XNOR2_X1 U499 ( .A(n516), .B(n442), .ZN(n490) );
  OR2_X1 U500 ( .A1(n742), .A2(n730), .ZN(n630) );
  XNOR2_X1 U501 ( .A(n553), .B(n554), .ZN(n680) );
  XNOR2_X1 U502 ( .A(n444), .B(n371), .ZN(n590) );
  NOR2_X1 U503 ( .A1(n570), .A2(n683), .ZN(n444) );
  INV_X1 U504 ( .A(n650), .ZN(n574) );
  XNOR2_X1 U505 ( .A(n549), .B(G475), .ZN(n436) );
  OR2_X1 U506 ( .A1(n715), .A2(G902), .ZN(n437) );
  INV_X1 U507 ( .A(KEYINPUT6), .ZN(n385) );
  BUF_X1 U508 ( .A(n665), .Z(n429) );
  XNOR2_X1 U509 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U510 ( .A(KEYINPUT122), .ZN(n463) );
  XNOR2_X1 U511 ( .A(n407), .B(n405), .ZN(n757) );
  XNOR2_X1 U512 ( .A(n406), .B(KEYINPUT111), .ZN(n405) );
  OR2_X1 U513 ( .A1(n680), .A2(n560), .ZN(n407) );
  INV_X1 U514 ( .A(KEYINPUT42), .ZN(n406) );
  XNOR2_X1 U515 ( .A(n616), .B(KEYINPUT79), .ZN(n447) );
  NOR2_X1 U516 ( .A1(n587), .A2(n570), .ZN(n571) );
  NOR2_X1 U517 ( .A1(n561), .A2(n560), .ZN(n648) );
  AND2_X1 U518 ( .A1(n398), .A2(n672), .ZN(n641) );
  XNOR2_X1 U519 ( .A(n711), .B(n710), .ZN(n712) );
  INV_X1 U520 ( .A(KEYINPUT53), .ZN(n426) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(n462) );
  NAND2_X1 U522 ( .A1(G210), .A2(n526), .ZN(n363) );
  OR2_X1 U523 ( .A1(n663), .A2(n662), .ZN(n364) );
  XOR2_X1 U524 ( .A(G472), .B(KEYINPUT72), .Z(n365) );
  XOR2_X1 U525 ( .A(n741), .B(n498), .Z(n366) );
  AND2_X1 U526 ( .A1(n416), .A2(n566), .ZN(n367) );
  XOR2_X1 U527 ( .A(n742), .B(KEYINPUT74), .Z(n368) );
  XOR2_X1 U528 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n369) );
  XNOR2_X1 U529 ( .A(KEYINPUT86), .B(KEYINPUT39), .ZN(n371) );
  XNOR2_X1 U530 ( .A(KEYINPUT89), .B(KEYINPUT0), .ZN(n372) );
  NOR2_X1 U531 ( .A1(n680), .A2(n682), .ZN(n373) );
  XOR2_X1 U532 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n374) );
  OR2_X1 U533 ( .A1(n629), .A2(n659), .ZN(n375) );
  XNOR2_X1 U534 ( .A(n517), .B(n516), .ZN(n520) );
  NOR2_X2 U535 ( .A1(n377), .A2(n376), .ZN(n627) );
  NAND2_X1 U536 ( .A1(n386), .A2(n626), .ZN(n376) );
  XNOR2_X2 U537 ( .A(n380), .B(n365), .ZN(n672) );
  NOR2_X1 U538 ( .A1(n582), .A2(n383), .ZN(n578) );
  XNOR2_X2 U539 ( .A(n459), .B(KEYINPUT88), .ZN(n383) );
  INV_X1 U540 ( .A(n384), .ZN(n533) );
  XNOR2_X2 U541 ( .A(n384), .B(n480), .ZN(n491) );
  AND2_X2 U542 ( .A1(n409), .A2(n454), .ZN(n453) );
  OR2_X2 U543 ( .A1(n701), .A2(n456), .ZN(n409) );
  XNOR2_X1 U544 ( .A(n733), .B(n392), .ZN(n701) );
  INV_X1 U545 ( .A(n672), .ZN(n622) );
  NAND2_X1 U546 ( .A1(n387), .A2(KEYINPUT44), .ZN(n386) );
  NAND2_X1 U547 ( .A1(n390), .A2(n753), .ZN(n387) );
  XNOR2_X2 U548 ( .A(n391), .B(n396), .ZN(n733) );
  XNOR2_X2 U549 ( .A(n524), .B(n394), .ZN(n391) );
  XNOR2_X1 U550 ( .A(n393), .B(n523), .ZN(n392) );
  XNOR2_X1 U551 ( .A(n396), .B(n395), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n621), .B(KEYINPUT100), .ZN(n398) );
  INV_X1 U553 ( .A(n400), .ZN(n602) );
  NAND2_X1 U554 ( .A1(n608), .A2(n400), .ZN(n610) );
  NOR2_X1 U555 ( .A1(n602), .A2(n399), .ZN(n621) );
  INV_X1 U556 ( .A(n620), .ZN(n399) );
  NAND2_X1 U557 ( .A1(n400), .A2(n676), .ZN(n624) );
  XNOR2_X1 U558 ( .A(n401), .B(n439), .ZN(n438) );
  NAND2_X1 U559 ( .A1(n440), .A2(n402), .ZN(n401) );
  XNOR2_X1 U560 ( .A(n559), .B(n374), .ZN(n402) );
  AND2_X1 U561 ( .A1(n409), .A2(n457), .ZN(n404) );
  NAND2_X1 U562 ( .A1(n408), .A2(n615), .ZN(n448) );
  NAND2_X1 U563 ( .A1(n408), .A2(n613), .ZN(n617) );
  XNOR2_X1 U564 ( .A(n410), .B(n369), .ZN(n519) );
  INV_X1 U565 ( .A(KEYINPUT44), .ZN(n414) );
  XNOR2_X2 U566 ( .A(n491), .B(n466), .ZN(n740) );
  NAND2_X1 U567 ( .A1(n453), .A2(n458), .ZN(n459) );
  XNOR2_X1 U568 ( .A(n415), .B(n490), .ZN(n477) );
  INV_X1 U569 ( .A(n524), .ZN(n415) );
  XNOR2_X1 U570 ( .A(n511), .B(n510), .ZN(n665) );
  XNOR2_X2 U571 ( .A(n419), .B(n475), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n451), .A2(n368), .ZN(n418) );
  NOR2_X2 U573 ( .A1(n602), .A2(n682), .ZN(n605) );
  NAND2_X1 U574 ( .A1(n757), .A2(n756), .ZN(n559) );
  NAND2_X1 U575 ( .A1(n438), .A2(n592), .ZN(n742) );
  NAND2_X1 U576 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U577 ( .A(n427), .B(n426), .ZN(G75) );
  NAND2_X1 U578 ( .A1(n462), .A2(n743), .ZN(n427) );
  XNOR2_X1 U579 ( .A(n584), .B(KEYINPUT1), .ZN(n600) );
  XNOR2_X2 U580 ( .A(n495), .B(n494), .ZN(n584) );
  XNOR2_X1 U581 ( .A(n430), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U582 ( .A1(n718), .A2(n726), .ZN(n430) );
  XNOR2_X1 U583 ( .A(n431), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U584 ( .A1(n706), .A2(n726), .ZN(n431) );
  NOR2_X2 U585 ( .A1(n730), .A2(n629), .ZN(n628) );
  XNOR2_X1 U586 ( .A(n485), .B(n484), .ZN(n632) );
  XNOR2_X1 U587 ( .A(n433), .B(n636), .ZN(G57) );
  NOR2_X2 U588 ( .A1(n635), .A2(n726), .ZN(n433) );
  NOR2_X1 U589 ( .A1(n619), .A2(n435), .ZN(n434) );
  INV_X1 U590 ( .A(n663), .ZN(n449) );
  XNOR2_X1 U591 ( .A(n628), .B(n452), .ZN(n451) );
  NAND2_X1 U592 ( .A1(n701), .A2(n363), .ZN(n458) );
  NAND2_X1 U593 ( .A1(n461), .A2(n606), .ZN(n460) );
  XNOR2_X1 U594 ( .A(n605), .B(n604), .ZN(n461) );
  XNOR2_X1 U595 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U596 ( .A(n717), .B(n716), .ZN(n718) );
  XOR2_X2 U597 ( .A(KEYINPUT4), .B(KEYINPUT66), .Z(n522) );
  XNOR2_X1 U598 ( .A(n709), .B(n468), .ZN(n710) );
  XOR2_X1 U599 ( .A(n708), .B(n707), .Z(n468) );
  INV_X1 U600 ( .A(n682), .ZN(n692) );
  INV_X1 U601 ( .A(n655), .ZN(n591) );
  INV_X1 U602 ( .A(KEYINPUT36), .ZN(n576) );
  NOR2_X1 U603 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U604 ( .A(n491), .B(n483), .ZN(n484) );
  XNOR2_X1 U605 ( .A(n576), .B(KEYINPUT87), .ZN(n577) );
  INV_X1 U606 ( .A(KEYINPUT59), .ZN(n714) );
  XNOR2_X1 U607 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U608 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n609) );
  XNOR2_X1 U609 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U610 ( .A(n366), .B(n505), .ZN(n724) );
  INV_X1 U611 ( .A(KEYINPUT32), .ZN(n616) );
  INV_X1 U612 ( .A(KEYINPUT63), .ZN(n636) );
  INV_X1 U613 ( .A(KEYINPUT40), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n469), .B(KEYINPUT14), .ZN(n470) );
  NAND2_X1 U615 ( .A1(G952), .A2(n470), .ZN(n698) );
  NOR2_X1 U616 ( .A1(G953), .A2(n698), .ZN(n595) );
  NAND2_X1 U617 ( .A1(n470), .A2(G902), .ZN(n471) );
  XOR2_X1 U618 ( .A(n471), .B(KEYINPUT93), .Z(n593) );
  OR2_X1 U619 ( .A1(n743), .A2(n593), .ZN(n472) );
  NOR2_X1 U620 ( .A1(G900), .A2(n472), .ZN(n473) );
  NOR2_X1 U621 ( .A1(n595), .A2(n473), .ZN(n556) );
  NAND2_X1 U622 ( .A1(G214), .A2(n526), .ZN(n474) );
  XNOR2_X1 U623 ( .A(KEYINPUT91), .B(n474), .ZN(n684) );
  NAND2_X1 U624 ( .A1(n540), .A2(G210), .ZN(n476) );
  XNOR2_X1 U625 ( .A(n477), .B(n476), .ZN(n485) );
  XNOR2_X1 U626 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U627 ( .A1(G227), .A2(n743), .ZN(n488) );
  XNOR2_X1 U628 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n493) );
  XNOR2_X1 U629 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U630 ( .A1(n743), .A2(G234), .ZN(n500) );
  XNOR2_X1 U631 ( .A(n500), .B(n499), .ZN(n534) );
  NAND2_X1 U632 ( .A1(G221), .A2(n534), .ZN(n504) );
  XOR2_X1 U633 ( .A(G110), .B(G119), .Z(n502) );
  XNOR2_X1 U634 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U635 ( .A(n504), .B(n503), .ZN(n505) );
  NOR2_X1 U636 ( .A1(G902), .A2(n724), .ZN(n511) );
  XOR2_X1 U637 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n508) );
  NAND2_X1 U638 ( .A1(n629), .A2(G234), .ZN(n506) );
  XNOR2_X1 U639 ( .A(n506), .B(KEYINPUT20), .ZN(n512) );
  NAND2_X1 U640 ( .A1(n512), .A2(G217), .ZN(n507) );
  XNOR2_X1 U641 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U642 ( .A(KEYINPUT98), .B(n509), .ZN(n510) );
  NAND2_X1 U643 ( .A1(G221), .A2(n512), .ZN(n513) );
  XOR2_X1 U644 ( .A(KEYINPUT21), .B(n513), .Z(n607) );
  INV_X1 U645 ( .A(n607), .ZN(n664) );
  NAND2_X1 U646 ( .A1(n584), .A2(n667), .ZN(n514) );
  XNOR2_X1 U647 ( .A(n514), .B(KEYINPUT99), .ZN(n620) );
  XOR2_X1 U648 ( .A(n522), .B(n521), .Z(n523) );
  INV_X1 U649 ( .A(n629), .ZN(n525) );
  XNOR2_X1 U650 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U651 ( .A(n529), .B(KEYINPUT7), .Z(n531) );
  XNOR2_X1 U652 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U653 ( .A(n533), .B(n532), .ZN(n536) );
  NAND2_X1 U654 ( .A1(G217), .A2(n534), .ZN(n535) );
  XNOR2_X1 U655 ( .A(n536), .B(n535), .ZN(n720) );
  NOR2_X1 U656 ( .A1(G902), .A2(n720), .ZN(n537) );
  XNOR2_X1 U657 ( .A(G478), .B(n537), .ZN(n564) );
  INV_X1 U658 ( .A(n564), .ZN(n567) );
  XNOR2_X1 U659 ( .A(n539), .B(n538), .ZN(n548) );
  NAND2_X1 U660 ( .A1(G214), .A2(n540), .ZN(n544) );
  XNOR2_X1 U661 ( .A(n542), .B(KEYINPUT12), .ZN(n543) );
  XNOR2_X1 U662 ( .A(n741), .B(KEYINPUT103), .ZN(n545) );
  XNOR2_X1 U663 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U664 ( .A(n548), .B(n547), .ZN(n715) );
  XNOR2_X1 U665 ( .A(KEYINPUT13), .B(KEYINPUT104), .ZN(n549) );
  NOR2_X1 U666 ( .A1(n590), .A2(n574), .ZN(n551) );
  XNOR2_X1 U667 ( .A(n552), .B(n551), .ZN(n756) );
  XOR2_X1 U668 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n554) );
  NOR2_X1 U669 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U670 ( .A1(n686), .A2(n688), .ZN(n553) );
  NAND2_X1 U671 ( .A1(n665), .A2(n607), .ZN(n555) );
  XNOR2_X1 U672 ( .A(n557), .B(KEYINPUT28), .ZN(n558) );
  NAND2_X1 U673 ( .A1(n558), .A2(n584), .ZN(n560) );
  INV_X1 U674 ( .A(n598), .ZN(n561) );
  INV_X1 U675 ( .A(KEYINPUT47), .ZN(n562) );
  NOR2_X1 U676 ( .A1(n648), .A2(n562), .ZN(n563) );
  NOR2_X1 U677 ( .A1(n564), .A2(n568), .ZN(n652) );
  INV_X1 U678 ( .A(n652), .ZN(n589) );
  NAND2_X1 U679 ( .A1(n574), .A2(n589), .ZN(n687) );
  INV_X1 U680 ( .A(n687), .ZN(n625) );
  NOR2_X1 U681 ( .A1(KEYINPUT47), .A2(n625), .ZN(n565) );
  NAND2_X1 U682 ( .A1(n648), .A2(n565), .ZN(n566) );
  NAND2_X1 U683 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U684 ( .A(n569), .B(KEYINPUT107), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n606), .A2(n571), .ZN(n572) );
  NAND2_X1 U686 ( .A1(n625), .A2(KEYINPUT47), .ZN(n573) );
  BUF_X1 U687 ( .A(n600), .Z(n668) );
  NAND2_X1 U688 ( .A1(n579), .A2(n668), .ZN(n580) );
  XNOR2_X1 U689 ( .A(n580), .B(KEYINPUT112), .ZN(n754) );
  NOR2_X1 U690 ( .A1(n684), .A2(n582), .ZN(n583) );
  XNOR2_X1 U691 ( .A(KEYINPUT108), .B(n583), .ZN(n585) );
  XOR2_X1 U692 ( .A(KEYINPUT1), .B(n584), .Z(n613) );
  NAND2_X1 U693 ( .A1(n585), .A2(n613), .ZN(n586) );
  XNOR2_X1 U694 ( .A(n586), .B(KEYINPUT43), .ZN(n588) );
  NAND2_X1 U695 ( .A1(n588), .A2(n587), .ZN(n657) );
  NOR2_X1 U696 ( .A1(n590), .A2(n589), .ZN(n655) );
  XOR2_X1 U697 ( .A(G898), .B(KEYINPUT92), .Z(n729) );
  NAND2_X1 U698 ( .A1(G953), .A2(n729), .ZN(n736) );
  NOR2_X1 U699 ( .A1(n593), .A2(n736), .ZN(n594) );
  NOR2_X1 U700 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U701 ( .A(KEYINPUT94), .B(n596), .Z(n597) );
  NAND2_X1 U702 ( .A1(n600), .A2(n667), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT34), .B(KEYINPUT78), .Z(n603) );
  XNOR2_X1 U704 ( .A(KEYINPUT71), .B(n603), .ZN(n604) );
  AND2_X1 U705 ( .A1(n607), .A2(n686), .ZN(n608) );
  NAND2_X1 U706 ( .A1(n429), .A2(n672), .ZN(n611) );
  NAND2_X1 U707 ( .A1(n429), .A2(n619), .ZN(n612) );
  NOR2_X1 U708 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U709 ( .A(KEYINPUT80), .B(n614), .ZN(n615) );
  NOR2_X1 U710 ( .A1(n429), .A2(n617), .ZN(n618) );
  NAND2_X1 U711 ( .A1(n619), .A2(n618), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n672), .A2(n623), .ZN(n676) );
  XNOR2_X1 U713 ( .A(KEYINPUT31), .B(n624), .ZN(n653) );
  AND2_X1 U714 ( .A1(n637), .A2(n370), .ZN(n626) );
  XNOR2_X2 U715 ( .A(n627), .B(KEYINPUT45), .ZN(n730) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n659) );
  NAND2_X1 U717 ( .A1(n713), .A2(G472), .ZN(n634) );
  XOR2_X1 U718 ( .A(KEYINPUT62), .B(KEYINPUT113), .Z(n631) );
  XNOR2_X1 U719 ( .A(G101), .B(n637), .ZN(G3) );
  XOR2_X1 U720 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n639) );
  NAND2_X1 U721 ( .A1(n356), .A2(n650), .ZN(n638) );
  XNOR2_X1 U722 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U723 ( .A(G104), .B(n640), .ZN(G6) );
  XOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U725 ( .A1(n356), .A2(n652), .ZN(n642) );
  XNOR2_X1 U726 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U727 ( .A(G107), .B(n644), .ZN(G9) );
  XOR2_X1 U728 ( .A(n645), .B(G110), .Z(G12) );
  XOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n652), .ZN(n646) );
  XNOR2_X1 U731 ( .A(n647), .B(n646), .ZN(G30) );
  NAND2_X1 U732 ( .A1(n648), .A2(n650), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n649), .B(G146), .ZN(G48) );
  NAND2_X1 U734 ( .A1(n653), .A2(n650), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n651), .B(n355), .ZN(G15) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n654), .B(G116), .ZN(G18) );
  XOR2_X1 U738 ( .A(G134), .B(n655), .Z(n656) );
  XNOR2_X1 U739 ( .A(KEYINPUT116), .B(n656), .ZN(G36) );
  XNOR2_X1 U740 ( .A(G140), .B(n657), .ZN(G42) );
  NAND2_X1 U741 ( .A1(n730), .A2(n659), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n658), .B(KEYINPUT84), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n742), .A2(n659), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U745 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n697) );
  NAND2_X1 U746 ( .A1(n429), .A2(n664), .ZN(n666) );
  XNOR2_X1 U747 ( .A(KEYINPUT49), .B(n666), .ZN(n674) );
  XNOR2_X1 U748 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U753 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U754 ( .A(n677), .B(KEYINPUT118), .Z(n678) );
  XNOR2_X1 U755 ( .A(KEYINPUT51), .B(n678), .ZN(n679) );
  NOR2_X1 U756 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U757 ( .A(n681), .B(KEYINPUT119), .ZN(n694) );
  NAND2_X1 U758 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U761 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(KEYINPUT120), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n713), .A2(G210), .ZN(n705) );
  BUF_X1 U768 ( .A(n701), .Z(n703) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n702) );
  NAND2_X1 U770 ( .A1(n722), .A2(G469), .ZN(n711) );
  XOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n708) );
  XNOR2_X1 U772 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n726), .A2(n712), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n713), .A2(G475), .ZN(n717) );
  NAND2_X1 U775 ( .A1(G478), .A2(n722), .ZN(n719) );
  NAND2_X1 U776 ( .A1(G217), .A2(n722), .ZN(n723) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n727) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(n727), .Z(n728) );
  NOR2_X1 U779 ( .A1(n729), .A2(n728), .ZN(n732) );
  NOR2_X1 U780 ( .A1(G953), .A2(n730), .ZN(n731) );
  NOR2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n739) );
  XOR2_X1 U782 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n735) );
  XNOR2_X1 U783 ( .A(n733), .B(G101), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n739), .B(n738), .ZN(G69) );
  XOR2_X1 U787 ( .A(n741), .B(n740), .Z(n745) );
  XNOR2_X1 U788 ( .A(n742), .B(n745), .ZN(n744) );
  NAND2_X1 U789 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U790 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U791 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U792 ( .A1(G953), .A2(n747), .ZN(n748) );
  NAND2_X1 U793 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U794 ( .A(KEYINPUT127), .B(n750), .Z(G72) );
  XOR2_X1 U795 ( .A(n751), .B(G122), .Z(G24) );
  XOR2_X1 U796 ( .A(G143), .B(n752), .Z(G45) );
  XNOR2_X1 U797 ( .A(G119), .B(n753), .ZN(G21) );
  XOR2_X1 U798 ( .A(n754), .B(G125), .Z(n755) );
  XNOR2_X1 U799 ( .A(KEYINPUT37), .B(n755), .ZN(G27) );
  XNOR2_X1 U800 ( .A(G131), .B(n756), .ZN(G33) );
  XNOR2_X1 U801 ( .A(G137), .B(n757), .ZN(G39) );
endmodule

