//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND3_X1   g034(.A1(new_n459), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n459), .B2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G101), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n459), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  AND3_X1   g047(.A1(new_n464), .A2(new_n466), .A3(G2105), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT67), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n464), .A2(new_n466), .A3(new_n459), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G124), .B1(G136), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n459), .B2(G114), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(G2104), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n475), .A2(G138), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(new_n490), .A3(new_n491), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(KEYINPUT71), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT72), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n515), .A2(new_n517), .A3(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n503), .A2(new_n516), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n519), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  AND3_X1   g103(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n515), .A2(new_n517), .A3(G543), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n518), .A2(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n505), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n535), .A2(G81), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n518), .A2(KEYINPUT9), .A3(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n531), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(new_n535), .B2(G91), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n537), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n555), .A2(new_n559), .A3(new_n562), .ZN(G299));
  OR2_X1    g138(.A1(new_n506), .A2(new_n512), .ZN(G303));
  OAI21_X1  g139(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n535), .A2(new_n568), .A3(G87), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT74), .B1(new_n523), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n518), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n501), .B2(new_n502), .ZN(new_n576));
  AND2_X1   g151(.A1(G73), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND4_X1   g155(.A1(G48), .A2(new_n508), .A3(new_n510), .A4(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n503), .A2(G86), .A3(new_n516), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n582), .B2(KEYINPUT77), .ZN(new_n583));
  OAI211_X1 g158(.A(KEYINPUT76), .B(G651), .C1(new_n576), .C2(new_n577), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n535), .A2(new_n585), .A3(G86), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n580), .A2(new_n583), .A3(new_n584), .A4(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n535), .A2(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G47), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n588), .B1(new_n589), .B2(new_n505), .C1(new_n537), .C2(new_n590), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT78), .Z(G290));
  NAND2_X1  g167(.A1(new_n535), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT10), .Z(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n531), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n518), .A2(G54), .B1(G651), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G284));
  OAI21_X1  g177(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n600), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g181(.A(new_n599), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n599), .A2(G559), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OR3_X1    g187(.A1(new_n612), .A2(KEYINPUT80), .A3(new_n600), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n612), .B2(new_n600), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G868), .C2(new_n548), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n474), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n475), .A2(G135), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  OR2_X1    g197(.A1(new_n460), .A2(new_n461), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n464), .A2(new_n466), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT13), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT15), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2435), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n635), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(G14), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT84), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n648), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n651), .B(new_n652), .C1(new_n646), .C2(new_n647), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n652), .A2(new_n645), .A3(new_n647), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  AOI22_X1  g243(.A1(new_n666), .A2(new_n667), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n663), .A2(new_n668), .A3(new_n665), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n669), .B(new_n670), .C1(new_n667), .C2(new_n666), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  INV_X1    g249(.A(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n673), .B(new_n677), .ZN(G229));
  XNOR2_X1  g253(.A(KEYINPUT86), .B(G16), .ZN(new_n679));
  MUX2_X1   g254(.A(G22), .B(G303), .S(new_n679), .Z(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G1971), .Z(new_n681));
  NOR2_X1   g256(.A1(G16), .A2(G23), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  MUX2_X1   g261(.A(G6), .B(G305), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n681), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT34), .Z(new_n691));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G25), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n474), .A2(G119), .B1(G131), .B2(new_n475), .ZN(new_n694));
  OR2_X1    g269(.A1(G95), .A2(G2105), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n693), .B1(new_n698), .B2(new_n692), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT35), .B(G1991), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n699), .B(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(new_n679), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT87), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n691), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n691), .A2(new_n708), .A3(new_n702), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n711));
  INV_X1    g286(.A(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(G29), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n480), .B2(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n713), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(KEYINPUT29), .ZN(new_n719));
  OAI21_X1  g294(.A(G2090), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G20), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n679), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT93), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT92), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT23), .Z(new_n725));
  NAND2_X1  g300(.A1(G299), .A2(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1956), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(KEYINPUT94), .B1(new_n720), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n719), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(new_n732), .A3(new_n717), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n548), .A2(new_n679), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G19), .B2(new_n679), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NOR2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n738), .A2(new_n739), .A3(G29), .ZN(new_n740));
  INV_X1    g315(.A(G160), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT30), .B(G28), .Z(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(G29), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G27), .A2(G29), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G164), .B2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2078), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n742), .A2(new_n743), .B1(new_n750), .B2(G11), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n746), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n692), .A2(G26), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT28), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n475), .A2(G140), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n756));
  NOR2_X1   g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n474), .B2(G128), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(new_n692), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT89), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n754), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(G2067), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(G2067), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n737), .B(new_n752), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n750), .B2(G11), .ZN(new_n769));
  NOR2_X1   g344(.A1(G4), .A2(G16), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n607), .B2(G16), .ZN(new_n771));
  MUX2_X1   g346(.A(G21), .B(G286), .S(G16), .Z(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(G1348), .B1(new_n772), .B2(G1966), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G1966), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G32), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n623), .A2(G105), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n475), .A2(G141), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G129), .B2(new_n474), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT27), .B(G1996), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n771), .A2(G1348), .B1(new_n735), .B2(new_n736), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n774), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n475), .A2(G139), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n624), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n459), .ZN(new_n791));
  MUX2_X1   g366(.A(G33), .B(new_n791), .S(G29), .Z(new_n792));
  AOI22_X1  g367(.A1(new_n792), .A2(G2072), .B1(new_n748), .B2(G2078), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n733), .A2(new_n769), .A3(new_n786), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n730), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G5), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G171), .B2(G16), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT90), .B(G1961), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n720), .A2(KEYINPUT94), .A3(new_n729), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n710), .A2(new_n795), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n792), .A2(G2072), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n621), .A2(new_n692), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(G311));
  AND3_X1   g379(.A1(new_n710), .A2(new_n795), .A3(new_n800), .ZN(new_n805));
  INV_X1    g380(.A(new_n802), .ZN(new_n806));
  INV_X1    g381(.A(new_n803), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n799), .ZN(G150));
  NAND2_X1  g383(.A1(new_n535), .A2(G93), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n809), .B1(new_n810), .B2(new_n505), .C1(new_n537), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G860), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n599), .A2(new_n608), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT38), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n548), .A2(new_n812), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n548), .A2(new_n812), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n816), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT95), .Z(new_n823));
  INV_X1    g398(.A(G860), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n814), .B1(new_n823), .B2(new_n825), .ZN(G145));
  XNOR2_X1  g401(.A(KEYINPUT98), .B(G37), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n791), .A2(KEYINPUT96), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n781), .B(new_n760), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(new_n497), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n497), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n791), .B(KEYINPUT96), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n474), .A2(G130), .B1(G142), .B2(new_n475), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n459), .A2(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n698), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n627), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT97), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n835), .A2(new_n841), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n621), .B(new_n741), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n480), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n827), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n846), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n835), .A2(new_n841), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT40), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G395));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n819), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n612), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n819), .B(KEYINPUT100), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n610), .B(KEYINPUT79), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n599), .B(G299), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(KEYINPUT41), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n860), .B2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT42), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n861), .A2(new_n862), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n859), .A2(new_n612), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n860), .A2(new_n863), .A3(new_n864), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G290), .B(G303), .ZN(new_n876));
  XNOR2_X1  g451(.A(G288), .B(G305), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n868), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n868), .B2(new_n875), .ZN(new_n881));
  OAI21_X1  g456(.A(G868), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n812), .A2(new_n600), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G295));
  NAND2_X1  g462(.A1(new_n882), .A2(new_n884), .ZN(G331));
  INV_X1    g463(.A(new_n827), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n819), .A2(G168), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n817), .A2(G286), .A3(new_n818), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G301), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(G171), .A3(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n866), .ZN(new_n896));
  INV_X1    g471(.A(new_n864), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n878), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n878), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n889), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n899), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(new_n900), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT43), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT43), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g489(.A(KEYINPUT103), .B(G1384), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n497), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n468), .A2(new_n471), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n760), .B(G2067), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT105), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n922), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n697), .A2(new_n700), .ZN(new_n929));
  INV_X1    g504(.A(G1996), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT104), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n781), .A2(new_n930), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n932), .A2(new_n781), .B1(new_n922), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n928), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G2067), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n760), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n923), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n928), .A2(new_n934), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n701), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n922), .B1(new_n940), .B2(new_n929), .ZN(new_n941));
  NOR3_X1   g516(.A1(G290), .A2(new_n923), .A3(G1986), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT48), .Z(new_n943));
  AND3_X1   g518(.A1(new_n939), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n932), .B(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n781), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n922), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT47), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT126), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n949), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n938), .B(new_n944), .C1(new_n951), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G8), .ZN(new_n957));
  NOR2_X1   g532(.A1(G166), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n959));
  NOR2_X1   g534(.A1(KEYINPUT107), .A2(KEYINPUT55), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n958), .B2(new_n959), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n497), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n497), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n732), .A3(new_n920), .A4(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n915), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n497), .B2(new_n963), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(new_n921), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n971), .B2(G1971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n962), .B1(new_n972), .B2(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n581), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n578), .A2(new_n974), .A3(new_n582), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G1981), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT49), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n978), .C1(G305), .C2(G1981), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G86), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n531), .A2(new_n511), .A3(new_n981), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n579), .A2(new_n578), .B1(new_n982), .B2(new_n585), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n983), .A2(new_n675), .A3(new_n584), .A4(new_n583), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n984), .B2(new_n976), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n920), .A2(new_n497), .A3(new_n963), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n986), .A2(KEYINPUT108), .A3(G8), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT108), .B1(new_n986), .B2(G8), .ZN(new_n988));
  OAI22_X1  g563(.A1(new_n980), .A2(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n683), .A2(G1976), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n990), .B(new_n992), .C1(new_n987), .C2(new_n988), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n986), .A2(G8), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(KEYINPUT108), .A3(G8), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n996), .A2(new_n997), .B1(G1976), .B2(new_n683), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n989), .B(new_n993), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n973), .B1(new_n1000), .B2(KEYINPUT110), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n972), .A2(G8), .A3(new_n962), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n964), .A2(new_n917), .ZN(new_n1003));
  INV_X1    g578(.A(G2078), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n915), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n920), .A4(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n965), .A2(new_n920), .A3(new_n967), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT119), .B(G1961), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT122), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n921), .B1(new_n1012), .B2(G2078), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(KEYINPUT122), .B2(new_n1004), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1013), .A2(new_n918), .A3(new_n1005), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1008), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G171), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n1006), .A2(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1003), .A2(KEYINPUT111), .A3(new_n920), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n970), .B2(new_n921), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1014), .A2(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(G301), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1018), .A2(new_n1026), .A3(KEYINPUT54), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n996), .A2(new_n997), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n990), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n989), .A4(new_n993), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1001), .A2(new_n1002), .A3(new_n1027), .A4(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n497), .A2(new_n966), .A3(new_n963), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n966), .B1(new_n497), .B2(new_n963), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n921), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT112), .A3(new_n743), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1009), .B2(G2084), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1040));
  INV_X1    g615(.A(G1966), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1037), .A2(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(new_n957), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1044), .B(KEYINPUT117), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1043), .A2(new_n1046), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1042), .A2(new_n957), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(new_n1049), .A3(KEYINPUT51), .A4(new_n1047), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1033), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1036), .A2(G1348), .B1(G2067), .B2(new_n986), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G299), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT57), .A4(new_n559), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1003), .A2(new_n920), .A3(new_n1005), .A4(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1060), .B(new_n1062), .C1(new_n1036), .C2(G1956), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1009), .A2(new_n728), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1065), .B2(new_n1062), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1056), .B1(new_n1067), .B2(KEYINPUT61), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1062), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1060), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1065), .A2(new_n1073), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT61), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1003), .A2(new_n930), .A3(new_n920), .A4(new_n1005), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n986), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1081), .A2(KEYINPUT116), .A3(new_n548), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1081), .A2(new_n548), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1086), .B2(KEYINPUT59), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1082), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1055), .A2(new_n607), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1055), .A2(new_n607), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1068), .A2(new_n1077), .A3(new_n1089), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1066), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1095), .B2(new_n1090), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1008), .A2(new_n1011), .A3(new_n1016), .A4(G301), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1019), .A2(new_n1103), .A3(G301), .A4(new_n1016), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g680(.A(KEYINPUT121), .B(G301), .C1(new_n1019), .C2(new_n1025), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1025), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(G171), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1100), .B1(new_n1110), .B2(KEYINPUT54), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT124), .B(new_n1112), .C1(new_n1113), .C2(new_n1105), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1054), .A2(new_n1099), .A3(new_n1111), .A4(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1043), .A2(G168), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1000), .A2(new_n973), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT63), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR4_X1   g694(.A1(new_n1042), .A2(KEYINPUT63), .A3(new_n957), .A4(G286), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(new_n1002), .A3(new_n1001), .A4(new_n1032), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n989), .A2(new_n991), .A3(new_n683), .ZN(new_n1122));
  INV_X1    g697(.A(new_n984), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1028), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND4_X1   g699(.A1(new_n1116), .A2(new_n1119), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1115), .A2(KEYINPUT125), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n1115), .B2(new_n1125), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1053), .A2(new_n1051), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1053), .A2(new_n1051), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1113), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1001), .A2(new_n1002), .A3(new_n1032), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1126), .A2(new_n1127), .A3(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(G290), .B(G1986), .Z(new_n1136));
  OAI211_X1 g711(.A(new_n939), .B(new_n941), .C1(new_n923), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n956), .B1(new_n1135), .B2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g713(.A1(G401), .A2(G227), .ZN(new_n1140));
  NAND2_X1  g714(.A1(new_n853), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g715(.A(G229), .ZN(new_n1142));
  OAI211_X1 g716(.A(G319), .B(new_n1142), .C1(new_n911), .C2(new_n912), .ZN(new_n1143));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1143), .ZN(G308));
  OR2_X1    g718(.A1(new_n911), .A2(new_n912), .ZN(new_n1145));
  INV_X1    g719(.A(new_n1140), .ZN(new_n1146));
  AOI21_X1  g720(.A(new_n1146), .B1(new_n847), .B2(new_n852), .ZN(new_n1147));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n1147), .A3(G319), .A4(new_n1142), .ZN(G225));
endmodule


