//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT11), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G134), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n191), .B2(G134), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(KEYINPUT64), .A3(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n187), .B1(new_n193), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n188), .A2(G137), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n191), .A2(G134), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n199), .A2(new_n200), .A3(new_n187), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n203), .B(G146), .C1(new_n204), .C2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT66), .A3(new_n207), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n198), .A2(new_n202), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(G146), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT0), .A4(G128), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT0), .B(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n210), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n187), .A2(KEYINPUT65), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n193), .B2(new_n197), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n188), .A2(KEYINPUT64), .A3(G137), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n188), .B2(G137), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n220), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n189), .A2(new_n192), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n219), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n214), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n208), .A2(new_n209), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n211), .A2(new_n215), .A3(new_n216), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n213), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(G131), .B1(new_n224), .B2(new_n226), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(new_n201), .ZN(new_n242));
  INV_X1    g056(.A(new_n219), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n193), .A2(new_n220), .A3(new_n197), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n225), .B1(new_n224), .B2(new_n226), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n237), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT28), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G237), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G210), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n249), .B(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n254), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n256), .B2(new_n258), .ZN(new_n261));
  OR2_X1    g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n242), .A2(new_n246), .A3(new_n237), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n248), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n214), .A2(new_n228), .A3(KEYINPUT30), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n242), .B2(new_n246), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n235), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n263), .ZN(new_n273));
  INV_X1    g087(.A(new_n262), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n266), .B2(new_n267), .ZN(new_n277));
  OAI21_X1  g091(.A(G472), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n272), .A2(new_n262), .A3(new_n263), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n272), .A2(new_n281), .A3(new_n262), .A4(new_n263), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n248), .A2(new_n265), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n274), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NOR2_X1   g100(.A1(G472), .A2(G902), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n278), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n278), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  INV_X1    g112(.A(G125), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(KEYINPUT72), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(G125), .A3(G140), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(KEYINPUT16), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT16), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n299), .B2(G140), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n206), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G125), .B(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n206), .ZN(new_n309));
  INV_X1    g123(.A(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G128), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n204), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n311), .B(new_n312), .C1(new_n314), .C2(KEYINPUT23), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(G110), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT24), .B(G110), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n313), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n311), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n307), .B(new_n309), .C1(new_n316), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n321), .A3(new_n317), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n315), .A2(G110), .ZN(new_n325));
  AND3_X1   g139(.A1(new_n303), .A2(new_n206), .A3(new_n305), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n306), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n323), .A2(new_n327), .A3(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n276), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n333), .A2(KEYINPUT25), .A3(new_n276), .A4(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G234), .ZN(new_n340));
  OAI21_X1  g154(.A(G217), .B1(new_n340), .B2(G902), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT70), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT73), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT73), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n345), .B(new_n342), .C1(new_n337), .C2(new_n338), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n333), .A2(new_n334), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n276), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n344), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G214), .B1(G237), .B2(G902), .ZN(new_n353));
  INV_X1    g167(.A(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n354), .B2(G107), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g170(.A(G107), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G104), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n355), .A2(new_n358), .A3(new_n362), .A4(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(G101), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n235), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G113), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n369));
  INV_X1    g183(.A(G116), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G119), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT79), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n229), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n372), .A2(new_n378), .B1(new_n229), .B2(new_n233), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n357), .A2(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n354), .A2(G107), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n363), .A2(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n379), .A2(KEYINPUT80), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT80), .B1(new_n379), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n367), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n367), .C1(new_n384), .C2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n205), .A2(KEYINPUT66), .A3(new_n207), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT66), .B1(new_n205), .B2(new_n207), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n211), .A2(new_n215), .A3(new_n216), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n299), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n219), .A2(G125), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n219), .A2(KEYINPUT81), .A3(G125), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT82), .B(G224), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n401), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n386), .A2(new_n405), .A3(new_n388), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n396), .A2(new_n397), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(new_n402), .B2(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n363), .A2(new_n382), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n379), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n387), .B(KEYINPUT8), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n372), .B1(new_n373), .B2(new_n230), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(new_n234), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n412), .B(new_n413), .C1(new_n415), .C2(new_n411), .ZN(new_n416));
  INV_X1    g230(.A(new_n409), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n396), .A2(new_n399), .A3(new_n400), .A4(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n410), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n390), .ZN(new_n420));
  OAI21_X1  g234(.A(G210), .B1(G237), .B2(G902), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n407), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n407), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n353), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n239), .A2(KEYINPUT76), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n205), .A2(new_n207), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT76), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n210), .A2(new_n429), .A3(new_n211), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n383), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n411), .B1(new_n212), .B2(new_n213), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT77), .B1(new_n244), .B2(new_n245), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT77), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n221), .A2(new_n437), .A3(new_n227), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n364), .A2(new_n243), .A3(new_n366), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n253), .A2(G227), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT74), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G140), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n431), .A2(new_n383), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n212), .A2(new_n213), .A3(new_n411), .ZN(new_n448));
  AOI221_X4 g262(.A(new_n446), .B1(new_n221), .B2(new_n227), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n221), .A2(new_n227), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT12), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n441), .B(new_n445), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n433), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n432), .B1(new_n240), .B2(new_n383), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n440), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n445), .B1(new_n458), .B2(new_n441), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n426), .B(new_n276), .C1(new_n454), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n441), .B1(new_n449), .B2(new_n452), .ZN(new_n461));
  INV_X1    g275(.A(new_n445), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n441), .A2(KEYINPUT78), .A3(new_n445), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT78), .B1(new_n441), .B2(new_n445), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(G469), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n426), .A2(new_n276), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G113), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n354), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT83), .B(G143), .ZN(new_n477));
  INV_X1    g291(.A(G214), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n478), .A2(G237), .A3(G953), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n203), .A2(KEYINPUT83), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n479), .A2(new_n481), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(new_n187), .C1(new_n479), .C2(new_n477), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT19), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n308), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n300), .A2(new_n302), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n488), .B(new_n206), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n486), .A2(new_n307), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n484), .B(KEYINPUT84), .C1(new_n479), .C2(new_n477), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n477), .A2(new_n479), .ZN(new_n495));
  INV_X1    g309(.A(new_n493), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(KEYINPUT84), .A3(new_n496), .A4(new_n484), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n300), .A2(G146), .A3(new_n302), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n494), .A2(new_n497), .B1(new_n309), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n476), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n483), .A2(new_n501), .A3(new_n485), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n326), .A2(new_n306), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT17), .B(G131), .C1(new_n480), .C2(new_n482), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n497), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n309), .A2(new_n498), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n508), .A3(new_n475), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(G475), .A2(G902), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT85), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n505), .A2(new_n508), .A3(new_n475), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n475), .B1(new_n505), .B2(new_n508), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n276), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT86), .B(G475), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n512), .A2(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n486), .A2(new_n307), .A3(new_n490), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n475), .B1(new_n508), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n511), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n511), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n370), .A2(G122), .ZN(new_n526));
  INV_X1    g340(.A(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(G116), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n528), .A3(new_n357), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT89), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT90), .B1(new_n526), .B2(KEYINPUT14), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT90), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n370), .A4(G122), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n528), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g352(.A(G128), .B(G143), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n188), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT13), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n204), .B2(G143), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n204), .A2(G143), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n203), .A2(KEYINPUT13), .A3(G128), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G134), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT88), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n357), .B1(new_n526), .B2(new_n528), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n529), .ZN(new_n552));
  INV_X1    g366(.A(new_n529), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT87), .B1(new_n553), .B2(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n188), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n541), .B1(new_n548), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G217), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n471), .A2(new_n558), .A3(G953), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n541), .B(new_n559), .C1(new_n548), .C2(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(G902), .B(new_n565), .C1(new_n561), .C2(new_n562), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g383(.A1(KEYINPUT91), .A2(G952), .ZN(new_n570));
  NAND2_X1  g384(.A1(KEYINPUT91), .A2(G952), .ZN(new_n571));
  AOI21_X1  g385(.A(G953), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n340), .B2(new_n252), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n573), .A2(KEYINPUT92), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(KEYINPUT92), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G898), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n253), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n276), .B1(G234), .B2(G237), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT93), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n576), .B(new_n585), .C1(new_n582), .C2(new_n580), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n518), .A2(new_n525), .A3(new_n569), .A4(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n425), .A2(new_n473), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n292), .A2(new_n297), .A3(new_n352), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n285), .A2(new_n276), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n593), .A2(G472), .B1(new_n285), .B2(new_n287), .ZN(new_n594));
  INV_X1    g408(.A(new_n472), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n596));
  INV_X1    g410(.A(new_n451), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n435), .B2(new_n440), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n462), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n599), .B2(new_n453), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n468), .B1(new_n600), .B2(new_n426), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n595), .B1(new_n601), .B2(new_n467), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(new_n352), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n594), .A2(KEYINPUT94), .A3(new_n352), .A4(new_n602), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n561), .A2(new_n562), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT33), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n561), .A2(new_n610), .A3(new_n562), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(G478), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n563), .A2(new_n564), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n564), .A2(new_n276), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n521), .A2(new_n522), .A3(new_n513), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n516), .A2(new_n517), .ZN(new_n619));
  INV_X1    g433(.A(new_n511), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n500), .B2(new_n509), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT20), .B1(new_n621), .B2(KEYINPUT85), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n521), .A2(new_n522), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n618), .B(new_n619), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n425), .A2(new_n625), .A3(new_n587), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n607), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n353), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n407), .A2(new_n420), .ZN(new_n631));
  INV_X1    g445(.A(new_n421), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n633), .B2(new_n422), .ZN(new_n634));
  INV_X1    g448(.A(new_n624), .ZN(new_n635));
  INV_X1    g449(.A(new_n569), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT95), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT95), .B1(new_n584), .B2(new_n586), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n607), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n339), .A2(new_n343), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n345), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n339), .A2(KEYINPUT73), .A3(new_n343), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n332), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n328), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n349), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n279), .A2(KEYINPUT31), .B1(new_n283), .B2(new_n274), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n652), .B2(new_n282), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n293), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n590), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT96), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G12));
  AND2_X1   g474(.A1(new_n292), .A2(new_n297), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n651), .A2(new_n473), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n582), .A2(G900), .A3(new_n253), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT97), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n576), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n637), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n661), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  XNOR2_X1  g483(.A(new_n665), .B(KEYINPUT39), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n602), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT99), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n633), .A2(new_n422), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n651), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n624), .A2(new_n636), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n630), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n274), .B1(new_n236), .B2(new_n247), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  INV_X1    g497(.A(new_n279), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n276), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n296), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n678), .A2(new_n681), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n673), .A2(new_n674), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT100), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NOR2_X1   g505(.A1(new_n625), .A2(new_n666), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n634), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n616), .B1(new_n518), .B2(new_n525), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n665), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT101), .B1(new_n696), .B2(new_n425), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n661), .A2(new_n662), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AOI21_X1  g514(.A(new_n595), .B1(new_n600), .B2(new_n426), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n600), .B2(new_n702), .ZN(new_n703));
  AOI211_X1 g517(.A(KEYINPUT102), .B(G902), .C1(new_n599), .C2(new_n453), .ZN(new_n704));
  OAI211_X1 g518(.A(KEYINPUT103), .B(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT10), .B1(new_n395), .B2(new_n411), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n243), .A2(new_n366), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n707), .A2(new_n433), .B1(new_n708), .B2(new_n364), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n441), .B1(new_n709), .B2(new_n597), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n462), .B1(new_n709), .B2(new_n439), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n240), .A2(new_n383), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n208), .B1(KEYINPUT76), .B2(new_n239), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n411), .B1(new_n713), .B2(new_n430), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n451), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n446), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n450), .A2(KEYINPUT12), .A3(new_n451), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n462), .A2(new_n710), .B1(new_n711), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT102), .B1(new_n719), .B2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n600), .A2(new_n702), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(G469), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT103), .B1(new_n722), .B2(new_n701), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n646), .A2(new_n647), .A3(new_n350), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n706), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n292), .A3(new_n297), .A4(new_n626), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT104), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n661), .A2(new_n728), .A3(new_n626), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n725), .A2(new_n641), .A3(new_n292), .A4(new_n297), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT105), .B(G116), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G18));
  OAI21_X1  g549(.A(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n634), .A3(new_n705), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n651), .A2(new_n589), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n292), .A3(new_n297), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NOR2_X1   g557(.A1(new_n706), .A2(new_n723), .ZN(new_n744));
  INV_X1    g558(.A(new_n640), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n624), .A2(new_n636), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n655), .A2(new_n746), .A3(new_n724), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n744), .A2(new_n747), .A3(new_n748), .A4(new_n634), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n640), .B(new_n569), .C1(new_n518), .C2(new_n525), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n594), .A2(new_n750), .A3(new_n352), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT106), .B1(new_n739), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NOR3_X1   g568(.A1(new_n696), .A2(new_n651), .A3(new_n655), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n740), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  NAND4_X1  g571(.A1(new_n633), .A2(new_n472), .A3(new_n353), .A4(new_n422), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n470), .A2(KEYINPUT107), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n601), .A2(new_n761), .A3(new_n467), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n352), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(KEYINPUT42), .A2(new_n617), .A3(new_n624), .A4(new_n665), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n290), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(new_n762), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n724), .A3(new_n758), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n292), .A3(new_n297), .A4(new_n692), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n770));
  AOI21_X1  g584(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n187), .ZN(G33));
  NAND2_X1  g586(.A1(new_n635), .A2(new_n636), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n666), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n292), .A3(new_n297), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  NOR2_X1   g590(.A1(new_n675), .A2(new_n630), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n635), .A2(new_n617), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n655), .A3(new_n679), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n778), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n426), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n787), .B2(new_n786), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n469), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n469), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n460), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n472), .A3(new_n670), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n785), .B(new_n796), .C1(new_n784), .C2(new_n783), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n472), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT47), .ZN(new_n800));
  INV_X1    g614(.A(new_n661), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n724), .A3(new_n692), .A4(new_n777), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NOR2_X1   g618(.A1(G952), .A2(G953), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT118), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n782), .A2(new_n577), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n744), .A2(new_n777), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n724), .B1(new_n296), .B2(new_n278), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT48), .ZN(new_n812));
  INV_X1    g626(.A(new_n572), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n686), .A2(new_n296), .A3(new_n352), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n808), .A2(new_n576), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(new_n815), .B2(new_n695), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n807), .A2(new_n724), .A3(new_n655), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n812), .B(new_n816), .C1(new_n739), .C2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n630), .A3(new_n677), .A4(new_n744), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT50), .Z(new_n821));
  NOR2_X1   g635(.A1(new_n617), .A2(new_n624), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n809), .A2(new_n656), .B1(new_n815), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n722), .A2(new_n460), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT110), .Z(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n800), .B1(new_n472), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n818), .A2(new_n778), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n819), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n828), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n820), .B(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n835), .A2(new_n836), .A3(new_n839), .A4(new_n823), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n834), .B1(new_n840), .B2(KEYINPUT51), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT117), .Z(new_n842));
  NOR3_X1   g656(.A1(new_n679), .A2(new_n595), .A3(new_n666), .ZN(new_n843));
  INV_X1    g657(.A(new_n767), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n425), .A2(new_n680), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n687), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n699), .A2(new_n668), .A3(new_n756), .A4(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n668), .A2(new_n699), .A3(new_n756), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT52), .A4(new_n846), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n353), .B(new_n745), .C1(new_n423), .C2(new_n424), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n773), .B2(new_n625), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n605), .A2(new_n606), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n591), .A3(new_n657), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n771), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n753), .A2(new_n733), .A3(new_n742), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n860), .A3(new_n730), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n569), .A2(new_n665), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n675), .A2(new_n630), .A3(new_n624), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n292), .A2(new_n297), .A3(new_n662), .A4(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n656), .A2(new_n844), .A3(new_n692), .A4(new_n759), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n775), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n775), .A2(new_n864), .A3(new_n868), .A4(new_n865), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT112), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n753), .A2(new_n733), .A3(new_n742), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n729), .B2(new_n727), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n869), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n859), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n871), .A2(new_n876), .ZN(new_n878));
  INV_X1    g692(.A(new_n848), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n854), .A2(new_n877), .B1(new_n880), .B2(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n875), .A4(new_n859), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n853), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n848), .B1(new_n871), .B2(new_n876), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n888), .A2(KEYINPUT114), .A3(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n882), .B1(new_n890), .B2(KEYINPUT54), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n806), .B1(new_n842), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n893));
  INV_X1    g707(.A(new_n814), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n678), .A2(new_n595), .A3(new_n630), .A4(new_n779), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n253), .A2(G952), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n890), .A2(G210), .A3(G902), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n391), .A2(new_n406), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n404), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  AND2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n853), .A2(new_n883), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT114), .B1(new_n888), .B2(KEYINPUT53), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n911), .B2(new_n276), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n890), .A2(KEYINPUT119), .A3(G902), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n632), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n899), .B(new_n906), .C1(new_n915), .C2(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(new_n890), .B(KEYINPUT54), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n468), .B(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n459), .B2(new_n454), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n789), .B(KEYINPUT120), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n899), .B1(new_n921), .B2(new_n923), .ZN(G54));
  AND2_X1   g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n913), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n510), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n510), .A2(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n912), .A2(new_n913), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT121), .ZN(new_n931));
  INV_X1    g745(.A(new_n899), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n912), .A2(new_n913), .A3(new_n933), .A4(new_n929), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT122), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n899), .B1(new_n926), .B2(new_n927), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n937), .A2(new_n938), .A3(new_n931), .A4(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(G60));
  AND2_X1   g754(.A1(new_n609), .A2(new_n611), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n614), .B(KEYINPUT59), .Z(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n891), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n899), .B(new_n944), .C1(new_n918), .C2(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n911), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n649), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n932), .C1(new_n347), .C2(new_n949), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT61), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n951), .B(new_n953), .ZN(G66));
  INV_X1    g768(.A(new_n858), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n873), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n253), .ZN(new_n957));
  INV_X1    g771(.A(new_n402), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n580), .B1(new_n958), .B2(new_n253), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n903), .B1(G898), .B2(new_n253), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  NOR2_X1   g778(.A1(new_n269), .A2(new_n271), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n488), .B1(new_n489), .B2(new_n487), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(G900), .B2(new_n253), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n690), .A2(new_n850), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n773), .A2(new_n625), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n777), .ZN(new_n973));
  OR4_X1    g787(.A1(new_n801), .A2(new_n724), .A3(new_n672), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n803), .A2(new_n797), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n970), .A2(new_n971), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT126), .B1(new_n977), .B2(new_n253), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n796), .A2(new_n845), .A3(new_n810), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT127), .Z(new_n980));
  INV_X1    g794(.A(new_n775), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n771), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n850), .A3(new_n976), .A4(new_n982), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n968), .B(new_n978), .C1(new_n253), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n253), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n967), .B1(new_n985), .B2(KEYINPUT126), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  OR3_X1    g802(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n988), .B1(new_n984), .B2(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G72));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n977), .B2(new_n956), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n274), .B1(new_n272), .B2(new_n263), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n993), .B1(new_n983), .B2(new_n956), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n273), .A2(new_n262), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n899), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n993), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n998), .A2(new_n995), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n881), .B2(new_n1002), .ZN(G57));
endmodule


