//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  INV_X1    g037(.A(G113), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(new_n470), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n466), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT67), .Z(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(KEYINPUT65), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n464), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT64), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(KEYINPUT3), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n480), .A2(new_n477), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n479), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n480), .A2(G2105), .A3(new_n488), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT66), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n493), .B2(G124), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT68), .Z(G162));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n477), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n486), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n477), .A2(G138), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n484), .A2(new_n485), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n484), .A2(KEYINPUT69), .A3(new_n485), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n461), .A2(new_n506), .A3(new_n500), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n499), .B1(new_n505), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n510), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g090(.A(G651), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT6), .B(G651), .Z(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n509), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n518), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n518), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT6), .B(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(G543), .A3(new_n533), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n524), .B1(new_n527), .B2(new_n528), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  AND3_X1   g111(.A1(new_n531), .A2(G543), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n526), .A2(G90), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  NAND2_X1  g119(.A1(new_n537), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n525), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n548), .A2(G651), .B1(new_n526), .B2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n525), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n537), .A2(G53), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n537), .B2(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(G299));
  XOR2_X1   g141(.A(new_n535), .B(KEYINPUT73), .Z(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n537), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n526), .A2(G87), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  AOI22_X1  g147(.A1(new_n509), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n518), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n509), .A2(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT74), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n540), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n526), .A2(G85), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  XNOR2_X1  g157(.A(KEYINPUT75), .B(G47), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n540), .B2(new_n582), .C1(new_n534), .C2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n527), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n525), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n588), .A2(new_n589), .B1(G651), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n534), .B2(KEYINPUT76), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(KEYINPUT76), .B2(new_n534), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n585), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n585), .B1(new_n598), .B2(G868), .ZN(G321));
  INV_X1    g175(.A(G286), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI211_X1 g178(.A(KEYINPUT77), .B(new_n603), .C1(new_n602), .C2(G299), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(KEYINPUT77), .B2(new_n603), .ZN(G297));
  XOR2_X1   g180(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n598), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n550), .A2(new_n602), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n597), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n493), .A2(G123), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n480), .A2(new_n477), .A3(new_n488), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G135), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n470), .A2(G2105), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n461), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n624), .A2(new_n625), .B1(new_n626), .B2(G2100), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n625), .B2(new_n624), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n626), .A2(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n620), .A2(new_n621), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT80), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT82), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n650), .A2(new_n651), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n655), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(KEYINPUT84), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  INV_X1    g247(.A(new_n669), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(KEYINPUT85), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n662), .A2(new_n663), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n669), .B2(new_n665), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n674), .B(new_n676), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n679), .B(new_n684), .ZN(G229));
  NOR2_X1   g260(.A1(G29), .A2(G35), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G162), .B2(G29), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT29), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(G2090), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G19), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n551), .B2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT92), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1341), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G21), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G168), .B2(new_n690), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT95), .B(G1966), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G5), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G171), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT96), .B(G1961), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n618), .A2(G29), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G28), .ZN(new_n705));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n704), .B2(G28), .ZN(new_n707));
  AND2_X1   g282(.A1(KEYINPUT31), .A2(G11), .ZN(new_n708));
  NOR2_X1   g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n705), .A2(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AOI21_X1  g286(.A(G29), .B1(new_n711), .B2(KEYINPUT24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(KEYINPUT24), .B2(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n474), .B2(new_n706), .ZN(new_n714));
  INV_X1    g289(.A(G2084), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n698), .A2(new_n702), .A3(new_n703), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n622), .A2(G105), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G141), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n489), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n493), .B2(G129), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n706), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n706), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G4), .A2(G16), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n598), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1348), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n694), .A2(new_n717), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n706), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n614), .A2(G140), .ZN(new_n736));
  OR2_X1    g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n493), .B2(G128), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(new_n706), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2067), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n690), .A2(G20), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT98), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT23), .ZN(new_n745));
  INV_X1    g320(.A(G299), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n690), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NOR2_X1   g323(.A1(G164), .A2(new_n706), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G27), .B2(new_n706), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n742), .A2(new_n748), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n706), .A2(G33), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  INV_X1    g332(.A(G139), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n489), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT93), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(new_n477), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n706), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G2072), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n727), .A2(new_n728), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n714), .A2(new_n715), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n733), .B(new_n754), .C1(KEYINPUT94), .C2(new_n770), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n689), .B(new_n771), .C1(KEYINPUT94), .C2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n688), .A2(G2090), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT97), .ZN(new_n774));
  INV_X1    g349(.A(G95), .ZN(new_n775));
  AND3_X1   g350(.A1(new_n775), .A2(new_n477), .A3(KEYINPUT87), .ZN(new_n776));
  AOI21_X1  g351(.A(KEYINPUT87), .B1(new_n775), .B2(new_n477), .ZN(new_n777));
  OAI221_X1 g352(.A(G2104), .B1(G107), .B2(new_n477), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G131), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n489), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n493), .B2(G119), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G29), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G25), .B2(G29), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT35), .B(G1991), .Z(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n690), .A2(G22), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n690), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n690), .A2(G23), .ZN(new_n797));
  INV_X1    g372(.A(G288), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n690), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT33), .B(G1976), .Z(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n690), .A2(G6), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n579), .B2(new_n690), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT90), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n799), .A2(new_n800), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n796), .A2(new_n801), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n810), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1986), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n790), .A2(new_n791), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT36), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n772), .A2(new_n774), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n819));
  XNOR2_X1  g394(.A(G150), .B(new_n819), .ZN(G311));
  NAND2_X1  g395(.A1(new_n526), .A2(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n534), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT101), .ZN(new_n824));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n525), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n540), .B1(new_n827), .B2(KEYINPUT100), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(KEYINPUT100), .B2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT104), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n598), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n550), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n550), .A2(new_n836), .A3(KEYINPUT103), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT103), .B1(new_n550), .B2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n830), .A2(new_n837), .A3(new_n839), .A4(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n835), .B(new_n844), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n833), .B1(new_n847), .B2(new_n849), .ZN(G145));
  INV_X1    g425(.A(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n477), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n489), .A2(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n493), .B2(G130), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n855), .A2(new_n624), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n624), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n785), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n785), .A2(new_n858), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n860), .A2(KEYINPUT105), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  INV_X1    g438(.A(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(new_n859), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n725), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n493), .A2(G128), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(new_n736), .A3(new_n738), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT69), .B1(new_n471), .B2(new_n500), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n507), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n499), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n740), .A2(G164), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n763), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n763), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n867), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n740), .A2(G164), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n764), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n725), .A3(new_n877), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n866), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n862), .A2(new_n865), .A3(new_n884), .A4(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(G162), .A2(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n494), .B(KEYINPUT68), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n474), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n619), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n891), .A3(new_n618), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n866), .B2(new_n885), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n885), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n880), .A2(KEYINPUT106), .A3(new_n884), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n899), .A2(new_n900), .A3(new_n860), .A4(new_n861), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n897), .A2(new_n901), .A3(KEYINPUT107), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT107), .B1(new_n897), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g480(.A1(new_n830), .A2(new_n602), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n844), .B(new_n610), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n598), .B(G299), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT108), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n908), .B(KEYINPUT41), .Z(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(G166), .B(new_n798), .ZN(new_n914));
  XNOR2_X1  g489(.A(G290), .B(new_n579), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n913), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n906), .B1(new_n918), .B2(new_n602), .ZN(G295));
  OAI21_X1  g494(.A(new_n906), .B1(new_n918), .B2(new_n602), .ZN(G331));
  NOR2_X1   g495(.A1(G168), .A2(G171), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n601), .B2(G171), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n844), .ZN(new_n923));
  NOR2_X1   g498(.A1(G286), .A2(G301), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n842), .B(new_n843), .C1(new_n924), .C2(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT109), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n922), .B2(new_n844), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n911), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n908), .A3(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n917), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n917), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n926), .A2(new_n909), .A3(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n923), .A2(new_n925), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n911), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n916), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n932), .A4(new_n931), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n932), .A3(new_n931), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n945), .B2(KEYINPUT43), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n934), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n946), .A2(KEYINPUT110), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT110), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G397));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G164), .B2(G1384), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT111), .B(G40), .Z(new_n953));
  OR2_X1    g528(.A1(new_n474), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n786), .A2(new_n789), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n786), .A2(new_n789), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n869), .A2(G2067), .ZN(new_n960));
  INV_X1    g535(.A(G2067), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n740), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n955), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT112), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n725), .B(G1996), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(G290), .B(G1986), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n959), .B(new_n967), .C1(new_n955), .C2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n474), .A2(new_n953), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n872), .B2(new_n873), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT116), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n874), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n715), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n979), .A2(new_n977), .A3(new_n715), .A4(new_n970), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT116), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(new_n952), .A3(new_n970), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n697), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n978), .A2(new_n981), .A3(G168), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G8), .ZN(new_n986));
  NOR2_X1   g561(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n985), .B(G8), .C1(KEYINPUT122), .C2(KEYINPUT51), .ZN(new_n989));
  NAND2_X1  g564(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n978), .A2(new_n981), .A3(new_n984), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(G8), .A3(new_n535), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(G166), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT55), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n970), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n1000));
  NOR3_X1   g575(.A1(G164), .A2(new_n951), .A3(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT113), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n982), .A2(new_n952), .A3(new_n1003), .A4(new_n970), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n795), .A3(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT114), .B1(new_n973), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n979), .A2(new_n977), .A3(new_n1009), .A4(new_n970), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n997), .B1(new_n1012), .B2(KEYINPUT115), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n999), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n579), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n997), .B1(new_n971), .B2(new_n970), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(G288), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1024), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(new_n1027), .C1(new_n1024), .C2(G288), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n973), .A2(new_n1006), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1008), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n997), .B1(new_n1005), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1032), .B2(new_n999), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT124), .B1(new_n1016), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1005), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1014), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n997), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1036), .B(new_n1033), .C1(new_n1039), .C2(new_n999), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G2078), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1042), .A2(KEYINPUT53), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1030), .A2(G1961), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n996), .A2(G171), .A3(new_n1041), .A4(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(G160), .A2(G40), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n952), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1051), .B2(new_n952), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n982), .B(new_n1047), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(new_n1044), .C1(new_n1042), .C2(KEYINPUT53), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G301), .B(KEYINPUT54), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1043), .A2(new_n1044), .A3(new_n1048), .A4(new_n1058), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n991), .A2(new_n993), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1067));
  XNOR2_X1  g642(.A(G299), .B(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n973), .B2(new_n1006), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT120), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n983), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1068), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n973), .B2(new_n1006), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n971), .A2(new_n970), .A3(new_n961), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1076), .B1(new_n597), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1045), .A2(new_n1073), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1067), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G299), .B(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n1070), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1076), .A2(new_n1086), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1080), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n598), .A3(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1076), .A2(KEYINPUT61), .A3(new_n1086), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1080), .A2(new_n1092), .A3(new_n598), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT58), .B(G1341), .Z(new_n1098));
  INV_X1    g673(.A(new_n971), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n954), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n983), .B2(G1996), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1101), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n551), .ZN(new_n1103));
  OR3_X1    g678(.A1(new_n1097), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1066), .B(new_n1087), .C1(new_n1096), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1097), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1107), .A2(new_n1090), .A3(new_n1095), .A4(new_n1094), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1066), .B1(new_n1108), .B2(new_n1087), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1062), .A2(new_n1035), .A3(KEYINPUT125), .A4(new_n1040), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1065), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(G1976), .B(G288), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1019), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1022), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1032), .A2(new_n999), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1029), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1032), .A2(new_n999), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n992), .A2(G8), .A3(new_n601), .ZN(new_n1119));
  AND4_X1   g694(.A1(KEYINPUT63), .A2(new_n1118), .A3(new_n1033), .A4(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1033), .B(new_n1119), .C1(new_n1039), .C2(new_n999), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n1123), .B2(KEYINPUT117), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1125), .A3(new_n1122), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1050), .B(new_n1112), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g704(.A(KEYINPUT118), .B(new_n1117), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n969), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n956), .A2(G1996), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT46), .Z(new_n1133));
  OAI21_X1  g708(.A(new_n955), .B1(new_n963), .B2(new_n867), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n967), .A2(new_n958), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n956), .B1(new_n1138), .B2(new_n962), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n967), .A2(new_n959), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n956), .A2(G1986), .A3(G290), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT48), .Z(new_n1142));
  AOI211_X1 g717(.A(new_n1137), .B(new_n1139), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1131), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g719(.A1(G401), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n942), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g721(.A(new_n1147), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1149));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1149), .ZN(G225));
endmodule


