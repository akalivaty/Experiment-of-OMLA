//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G236), .A4(G238), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G101), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n463), .A2(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n464), .A2(new_n472), .A3(new_n465), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT71), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(new_n476), .A3(G125), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n473), .A2(new_n476), .A3(KEYINPUT72), .A4(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT70), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n471), .B1(new_n482), .B2(new_n485), .ZN(G160));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT73), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n466), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n466), .A2(new_n469), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g067(.A1(G124), .A2(new_n490), .B1(new_n492), .B2(G136), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n488), .A2(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n460), .A2(new_n461), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n476), .A3(new_n473), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n483), .A2(KEYINPUT4), .A3(G138), .A4(new_n484), .ZN(new_n500));
  NAND2_X1  g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n466), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(new_n469), .B2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n499), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT74), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G62), .A3(G651), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n515), .A2(new_n516), .A3(new_n521), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n515), .A2(KEYINPUT75), .A3(G543), .A4(new_n516), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(G51), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT7), .Z(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n524), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(KEYINPUT76), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n523), .A2(G89), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n532), .A2(new_n542), .A3(new_n543), .A4(new_n538), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n511), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT77), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n524), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n530), .A2(new_n531), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n552), .A2(G52), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  NAND2_X1  g129(.A1(new_n523), .A2(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT5), .B(G543), .Z(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT78), .B1(new_n559), .B2(G651), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n521), .A2(G56), .ZN(new_n562));
  AOI211_X1 g137(.A(new_n561), .B(new_n511), .C1(new_n562), .C2(new_n556), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n555), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n530), .A2(G43), .A3(new_n531), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND4_X1  g146(.A1(new_n517), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n523), .A2(G91), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n528), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n572), .A2(new_n574), .A3(new_n575), .A4(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  AND2_X1   g155(.A1(new_n541), .A2(new_n544), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND3_X1  g157(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n523), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n517), .A2(KEYINPUT79), .A3(G48), .A4(G543), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(new_n590), .B1(G86), .B2(new_n523), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n511), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n552), .A2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n557), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n523), .A2(G85), .B1(new_n599), .B2(G651), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(G290));
  NAND3_X1  g176(.A1(G301), .A2(KEYINPUT80), .A3(G868), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(G171), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n523), .A2(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n530), .A2(G54), .A3(new_n531), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(new_n511), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n610), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n602), .B(new_n605), .C1(G868), .C2(new_n616), .ZN(G284));
  OAI211_X1 g192(.A(new_n602), .B(new_n605), .C1(G868), .C2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(KEYINPUT81), .B1(new_n604), .B2(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(KEYINPUT81), .B2(new_n619), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(KEYINPUT81), .B2(new_n619), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n564), .A2(new_n565), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n626), .A2(new_n627), .B1(new_n604), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n627), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n473), .A2(new_n476), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(new_n470), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  AOI22_X1  g213(.A1(G123), .A2(new_n490), .B1(new_n492), .B2(G135), .ZN(new_n639));
  OAI221_X1 g214(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(G156));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT83), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT17), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n667), .B2(new_n663), .ZN(new_n668));
  INV_X1    g243(.A(new_n661), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n663), .A3(new_n661), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n642), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2100), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G26), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  AOI22_X1  g271(.A1(G128), .A2(new_n490), .B1(new_n492), .B2(G140), .ZN(new_n697));
  OAI221_X1 g272(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n699), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G2067), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G28), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n703), .B2(KEYINPUT30), .ZN(new_n705));
  OR2_X1    g280(.A1(KEYINPUT31), .A2(G11), .ZN(new_n706));
  NAND2_X1  g281(.A1(KEYINPUT31), .A2(G11), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n641), .B2(new_n694), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G164), .A2(new_n694), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G27), .B2(new_n694), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT93), .B(G2078), .Z(new_n713));
  OAI21_X1  g288(.A(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n694), .A2(G33), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT25), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G139), .B2(new_n492), .ZN(new_n718));
  NAND2_X1  g293(.A1(G115), .A2(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G127), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n632), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(new_n485), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n715), .B1(new_n724), .B2(new_n694), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n694), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n694), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT29), .B(G2090), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n725), .A2(G2072), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n712), .A2(new_n713), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n726), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NOR2_X1   g310(.A1(G171), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G5), .B2(new_n735), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n714), .B(new_n733), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n735), .A2(G4), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n616), .B2(new_n735), .ZN(new_n744));
  INV_X1    g319(.A(G1348), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n735), .A2(G19), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n566), .B2(new_n735), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n694), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n749), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n738), .A2(new_n742), .A3(new_n746), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n737), .A2(new_n734), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n735), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n735), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n760), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n755), .A2(G2084), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT86), .Z(new_n768));
  NOR3_X1   g343(.A1(new_n758), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G105), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(new_n470), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n772), .A2(new_n469), .A3(G105), .A4(G2104), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G141), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n491), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G129), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n489), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n776), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n776), .B2(new_n781), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT90), .Z(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G29), .B2(G32), .ZN(new_n789));
  INV_X1    g364(.A(G1996), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT91), .B(KEYINPUT27), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n769), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n735), .A2(G6), .ZN(new_n796));
  INV_X1    g371(.A(G305), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n735), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n735), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n735), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n735), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n735), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT33), .B(G1976), .Z(new_n806));
  AOI22_X1  g381(.A1(new_n802), .A2(G1971), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n807), .B(new_n808), .C1(G1971), .C2(new_n802), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n800), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT85), .Z(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n810), .B(KEYINPUT85), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G24), .ZN(new_n816));
  INV_X1    g391(.A(G290), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n818), .A2(G1986), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(G1986), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n694), .A2(G25), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n490), .A2(G119), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n492), .A2(G131), .ZN(new_n823));
  OAI221_X1 g398(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n821), .B1(new_n826), .B2(new_n694), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT35), .B(G1991), .Z(new_n828));
  XOR2_X1   g403(.A(new_n827), .B(new_n828), .Z(new_n829));
  NOR3_X1   g404(.A1(new_n819), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n813), .A2(new_n815), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n813), .A2(new_n815), .A3(new_n833), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n795), .B1(new_n832), .B2(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n793), .A2(new_n794), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n769), .ZN(G150));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n557), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n511), .B1(new_n841), .B2(KEYINPUT94), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(new_n839), .C1(new_n557), .C2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n530), .A2(G55), .A3(new_n531), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n523), .A2(G93), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n842), .A2(new_n844), .B1(G93), .B2(new_n523), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n846), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n566), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n848), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n616), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n859), .A2(new_n860), .A3(G860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n849), .A2(new_n852), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n861), .A2(new_n864), .ZN(G145));
  NOR2_X1   g440(.A1(new_n462), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n866), .A2(new_n867), .B1(new_n491), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n489), .A2(KEYINPUT96), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT96), .B1(new_n489), .B2(new_n870), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n634), .B(new_n873), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n786), .A2(new_n724), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n723), .A2(new_n785), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n699), .B(new_n508), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n826), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n875), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n881), .ZN(new_n884));
  INV_X1    g459(.A(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n878), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G160), .B(new_n641), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G162), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n883), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(KEYINPUT97), .A3(new_n892), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g473(.A1(new_n862), .A2(new_n604), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n855), .B(new_n625), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n572), .A2(new_n578), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n574), .A2(new_n575), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n615), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n613), .B1(new_n608), .B2(new_n609), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(G299), .A3(new_n611), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n904), .A2(G299), .A3(new_n611), .ZN(new_n910));
  AOI21_X1  g485(.A(G299), .B1(new_n904), .B2(new_n611), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n908), .A2(KEYINPUT98), .B1(new_n900), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT98), .B2(new_n908), .ZN(new_n916));
  XNOR2_X1  g491(.A(G305), .B(G290), .ZN(new_n917));
  XNOR2_X1  g492(.A(G166), .B(G288), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT42), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n916), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n899), .B1(new_n921), .B2(new_n604), .ZN(G295));
  OAI21_X1  g497(.A(new_n899), .B1(new_n921), .B2(new_n604), .ZN(G331));
  NOR3_X1   g498(.A1(new_n853), .A2(new_n854), .A3(G286), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n848), .A2(KEYINPUT95), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n851), .B1(new_n850), .B2(new_n846), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n628), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n566), .A2(new_n846), .A3(new_n850), .ZN(new_n928));
  AOI21_X1  g503(.A(G168), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(G301), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(G286), .B1(new_n853), .B2(new_n854), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(G168), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(G171), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n906), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT101), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n906), .A2(new_n936), .A3(new_n909), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n930), .B2(new_n933), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT102), .B(new_n938), .C1(new_n930), .C2(new_n933), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n919), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n931), .A2(new_n932), .A3(G171), .ZN(new_n944));
  AOI21_X1  g519(.A(G171), .B1(new_n931), .B2(new_n932), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n914), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n919), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n934), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G37), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT103), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n943), .A2(new_n950), .A3(new_n954), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n934), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n919), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n951), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n943), .A2(new_n950), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  OAI221_X1 g540(.A(KEYINPUT44), .B1(new_n959), .B2(new_n958), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n508), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT45), .B1(new_n969), .B2(KEYINPUT104), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(KEYINPUT104), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n482), .A2(new_n485), .ZN(new_n972));
  OAI221_X1 g547(.A(G40), .B1(new_n468), .B2(new_n470), .C1(new_n463), .C2(new_n467), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT105), .Z(new_n977));
  INV_X1    g552(.A(G1986), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n817), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT106), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT48), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n699), .A2(G2067), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(G1996), .B2(new_n785), .ZN(new_n986));
  INV_X1    g561(.A(new_n786), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(G1996), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n825), .B(new_n828), .Z(new_n989));
  OAI21_X1  g564(.A(new_n977), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n977), .A2(KEYINPUT48), .A3(new_n980), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n982), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n826), .A2(new_n828), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n984), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n977), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n977), .A2(new_n790), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n985), .A2(new_n785), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n996), .A2(new_n997), .B1(new_n977), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n997), .B2(new_n996), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n992), .B(new_n995), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n589), .A2(new_n590), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n523), .A2(G86), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n593), .B1(new_n1006), .B2(KEYINPUT113), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n591), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n691), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT112), .B(G1981), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n797), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1013), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1010), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n973), .B1(new_n482), .B2(new_n485), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n506), .B1(new_n497), .B2(new_n498), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n1019), .B2(new_n503), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1022), .A2(KEYINPUT111), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1021), .B2(G8), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1014), .A2(new_n1017), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n804), .A2(G1976), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1028), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G166), .A2(new_n1023), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT55), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(KEYINPUT109), .A3(KEYINPUT55), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT110), .B1(new_n1036), .B2(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1042), .B(new_n1043), .C1(G166), .C2(new_n1023), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1018), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1020), .A2(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT108), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n969), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(new_n1046), .A4(new_n1018), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1020), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1018), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1054), .A2(G1971), .B1(G2090), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1045), .A2(new_n1059), .A3(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1035), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1028), .A2(new_n1030), .A3(new_n804), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1013), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1027), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1028), .A2(new_n1060), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1023), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1045), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1055), .A2(new_n1057), .A3(new_n750), .A4(new_n1018), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT115), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT50), .B(G1384), .C1(new_n1019), .C2(new_n503), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1056), .B1(new_n508), .B2(new_n968), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n750), .A4(new_n1018), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1051), .A2(new_n1046), .A3(new_n1018), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n763), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT63), .B1(new_n1070), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1059), .A2(G8), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT63), .B(new_n1081), .C1(new_n1083), .C2(new_n1045), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1065), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1064), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n901), .B(new_n902), .C1(KEYINPUT116), .C2(KEYINPUT57), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n572), .A2(KEYINPUT116), .A3(new_n578), .ZN(new_n1089));
  NAND3_X1  g664(.A1(G299), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1058), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1051), .A2(new_n1046), .A3(new_n1018), .A4(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n745), .A2(new_n1058), .B1(new_n1022), .B2(new_n701), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n615), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1094), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1058), .A2(new_n745), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1022), .A2(new_n701), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT60), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n1108), .B2(new_n615), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n616), .C1(new_n1101), .C2(KEYINPUT60), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT58), .B(G1341), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1078), .A2(G1996), .B1(new_n1022), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n566), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT59), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1103), .A2(KEYINPUT61), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1100), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1956), .B1(new_n1075), .B2(new_n1018), .ZN(new_n1122));
  AND4_X1   g697(.A1(new_n1051), .A2(new_n1046), .A3(new_n1018), .A4(new_n1096), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1092), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1103), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1128), .B(KEYINPUT61), .C1(new_n1124), .C2(new_n1103), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1119), .B(new_n1121), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1105), .B1(new_n1115), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  AOI21_X1  g707(.A(G1961), .B1(new_n1075), .B2(new_n1018), .ZN(new_n1133));
  INV_X1    g708(.A(G2078), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1135), .A2(new_n1048), .A3(new_n975), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT122), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1135), .A2(new_n975), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1051), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1058), .A2(new_n734), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1054), .A2(new_n1134), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1137), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1132), .B1(new_n1145), .B2(G301), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1142), .A2(new_n1137), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n971), .A2(new_n1138), .B1(new_n1058), .B2(new_n734), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1148), .A2(G301), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1146), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1080), .A2(KEYINPUT120), .ZN(new_n1156));
  AOI22_X1  g731(.A1(KEYINPUT115), .A2(new_n1071), .B1(new_n1078), .B2(new_n763), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n1077), .ZN(new_n1159));
  AOI21_X1  g734(.A(G286), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1023), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G168), .A2(new_n1023), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1156), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1164), .B(G8), .C1(new_n1080), .C2(G286), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1145), .B2(G301), .ZN(new_n1168));
  AOI21_X1  g743(.A(G2078), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1151), .B1(new_n1169), .B2(KEYINPUT53), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1151), .B(KEYINPUT125), .C1(new_n1169), .C2(KEYINPUT53), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1172), .A2(G171), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1161), .A2(new_n1166), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1131), .A2(new_n1155), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n1161), .B2(new_n1166), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1161), .A2(new_n1166), .A3(new_n1177), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1158), .B1(new_n1157), .B2(new_n1077), .ZN(new_n1182));
  AND4_X1   g757(.A1(new_n1158), .A2(new_n1072), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1183));
  OAI21_X1  g758(.A(G168), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1164), .B1(new_n1184), .B2(G8), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1179), .B(KEYINPUT62), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1176), .B1(new_n1181), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1070), .B(KEYINPUT124), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1086), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n817), .A2(new_n978), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n977), .B1(new_n980), .B2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g769(.A(new_n1194), .B(KEYINPUT107), .Z(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n990), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1003), .B1(new_n1192), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g772(.A1(G227), .A2(new_n458), .ZN(new_n1199));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1200));
  OR2_X1    g774(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g777(.A1(G229), .A2(G401), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g779(.A1(new_n961), .A2(new_n1205), .A3(new_n897), .ZN(G308));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n1205), .A3(new_n897), .ZN(G225));
endmodule


