//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  OAI21_X1  g007(.A(G128), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n187), .A3(new_n191), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n189), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(new_n191), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n194), .A2(new_n197), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT3), .A2(G107), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT74), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G104), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT74), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT3), .A2(G107), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(G104), .B2(new_n204), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(G104), .A2(G107), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT74), .B(G104), .ZN(new_n216));
  OAI211_X1 g030(.A(G101), .B(new_n215), .C1(new_n216), .C2(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n203), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n201), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n196), .A2(KEYINPUT76), .A3(KEYINPUT1), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT64), .A2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT64), .A2(G146), .ZN(new_n225));
  OAI21_X1  g039(.A(G143), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n198), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n222), .A2(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n202), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n214), .B(new_n217), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n233), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n237), .A2(new_n239), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n236), .B1(new_n243), .B2(G137), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(G137), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n244), .A2(new_n241), .A3(new_n240), .A4(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n238), .A3(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n232), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT12), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n232), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT12), .B1(new_n232), .B2(new_n248), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n242), .A2(new_n247), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n250), .B(new_n256), .C1(new_n219), .C2(new_n231), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT81), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n211), .A2(KEYINPUT75), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n208), .A2(KEYINPUT74), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n206), .A2(G104), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n204), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g077(.A(G107), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G104), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT3), .A2(G107), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(KEYINPUT4), .B(new_n259), .C1(new_n262), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n262), .A2(new_n267), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n211), .ZN(new_n271));
  INV_X1    g085(.A(new_n259), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n201), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n226), .A2(new_n227), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n226), .A2(new_n279), .A3(new_n227), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(new_n201), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n276), .B1(new_n195), .B2(new_n196), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n278), .A2(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT10), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n274), .A2(new_n283), .B1(new_n231), .B2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n214), .A2(new_n217), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT77), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n201), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n288));
  INV_X1    g102(.A(new_n196), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n224), .A2(new_n225), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n187), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n229), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT10), .A4(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n214), .A2(KEYINPUT10), .A3(new_n217), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT77), .B1(new_n203), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n285), .A2(new_n296), .A3(new_n256), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G140), .ZN(new_n298));
  INV_X1    g112(.A(G227), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G953), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n298), .B(new_n300), .Z(new_n301));
  NAND4_X1  g115(.A1(new_n254), .A2(new_n258), .A3(new_n297), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n301), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n285), .A2(new_n296), .A3(new_n256), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n256), .B1(new_n285), .B2(new_n296), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT80), .B(G469), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n255), .A2(new_n257), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n304), .ZN(new_n315));
  INV_X1    g129(.A(new_n305), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n297), .A3(new_n301), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n308), .A3(new_n321), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n322), .A2(KEYINPUT79), .A3(G469), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT79), .B1(new_n322), .B2(G469), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n311), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G217), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(G234), .B2(new_n308), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT71), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT16), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(new_n329), .A3(KEYINPUT71), .A4(G125), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n333), .C1(new_n332), .C2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n189), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n201), .A2(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G128), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G110), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n339), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT24), .B(G110), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n337), .A2(new_n189), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n349), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n346), .B2(G110), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n199), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G953), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G221), .A3(G234), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT72), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT22), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n361), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n233), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n367), .A3(G137), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n359), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n351), .A3(new_n358), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n375), .B2(new_n308), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n377), .B(G902), .C1(new_n372), .C2(new_n374), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n327), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n375), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n327), .A2(G902), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(G472), .A2(G902), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT31), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n278), .A2(new_n280), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n282), .A2(new_n281), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n248), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n342), .A2(G116), .ZN(new_n389));
  INV_X1    g203(.A(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G119), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT2), .B(G113), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n246), .A2(G131), .ZN(new_n396));
  INV_X1    g210(.A(G131), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n235), .B2(new_n245), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n292), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT68), .B1(new_n396), .B2(new_n398), .ZN(new_n404));
  INV_X1    g218(.A(new_n398), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT68), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n405), .B(new_n406), .C1(new_n246), .C2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n292), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT30), .B1(new_n408), .B2(new_n388), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n410), .B2(new_n394), .ZN(new_n411));
  INV_X1    g225(.A(G237), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n360), .A3(G210), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT27), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT26), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n211), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n385), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n408), .A2(new_n388), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n394), .A3(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(new_n385), .A3(new_n401), .A4(new_n416), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n401), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n394), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n388), .A2(KEYINPUT28), .A3(new_n400), .A4(new_n395), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT32), .B(new_n384), .C1(new_n417), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n422), .A2(new_n401), .A3(new_n416), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT31), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n423), .A3(new_n430), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT32), .B1(new_n436), .B2(new_n384), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n395), .B1(new_n388), .B2(new_n400), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n402), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT69), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(KEYINPUT28), .C1(new_n402), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n425), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n444), .A2(new_n445), .A3(new_n429), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n411), .A2(new_n416), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n428), .B2(new_n429), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n308), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G472), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n383), .B1(new_n438), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT9), .B(G234), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G221), .B1(new_n453), .B2(G902), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n325), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n265), .B(new_n266), .C1(new_n216), .C2(new_n204), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n214), .A2(KEYINPUT4), .B1(new_n456), .B2(new_n259), .ZN(new_n457));
  INV_X1    g271(.A(new_n268), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n394), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n460), .B(G113), .C1(KEYINPUT5), .C2(new_n389), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n392), .A2(new_n393), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n286), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n214), .A2(new_n461), .A3(new_n462), .A4(new_n217), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT83), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(KEYINPUT84), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n459), .A2(new_n469), .A3(new_n465), .A4(new_n467), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n468), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n386), .A2(G125), .A3(new_n387), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n292), .A2(new_n334), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n360), .A2(G224), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n469), .B(KEYINPUT8), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n461), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n218), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n485), .B2(new_n466), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(KEYINPUT7), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n479), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n479), .B2(new_n488), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n477), .A2(KEYINPUT85), .A3(new_n478), .A4(new_n487), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n474), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n493), .A2(new_n308), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n482), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n496), .A3(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G214), .B1(G237), .B2(G902), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n338), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n412), .A2(new_n360), .A3(G214), .ZN(new_n506));
  NOR2_X1   g320(.A1(KEYINPUT86), .A2(G143), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n397), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n337), .A2(new_n189), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n353), .A2(KEYINPUT90), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT17), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n505), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n208), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n336), .A2(KEYINPUT87), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT87), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n356), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G146), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n524), .A2(new_n357), .B1(new_n509), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n516), .A2(KEYINPUT18), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n520), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT19), .B1(new_n521), .B2(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT88), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n336), .A2(KEYINPUT19), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(KEYINPUT19), .C1(new_n521), .C2(new_n523), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n532), .A2(new_n199), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n352), .B1(new_n510), .B2(new_n512), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n536), .A2(new_n537), .B1(new_n526), .B2(new_n527), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n530), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n537), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n541), .A2(new_n539), .A3(new_n528), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n529), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G475), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n308), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n529), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n520), .B1(new_n518), .B2(new_n528), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n308), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G475), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n544), .A4(new_n308), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n360), .A2(G952), .ZN(new_n554));
  NAND2_X1  g368(.A1(G234), .A2(G237), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT95), .Z(new_n557));
  XOR2_X1   g371(.A(KEYINPUT21), .B(G898), .Z(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(G902), .A3(G953), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n201), .B2(G143), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n187), .A2(KEYINPUT13), .A3(G128), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n569), .B(new_n570), .C1(G128), .C2(new_n187), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G134), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  XNOR2_X1  g387(.A(G128), .B(G143), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n243), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n576), .A3(G134), .ZN(new_n577));
  XNOR2_X1  g391(.A(G116), .B(G122), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n264), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n573), .A2(new_n575), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G122), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G116), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n264), .B1(new_n582), .B2(KEYINPUT14), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n578), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n574), .B(new_n243), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n584), .A2(KEYINPUT92), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT92), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n453), .A2(new_n326), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n580), .B(new_n589), .C1(new_n586), .C2(new_n587), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT93), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n595), .B(G902), .C1(new_n591), .C2(new_n592), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n567), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n567), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n553), .A2(new_n561), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n503), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n455), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  INV_X1    g418(.A(new_n454), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n322), .A2(G469), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n322), .A2(KEYINPUT79), .A3(G469), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n605), .B1(new_n610), .B2(new_n311), .ZN(new_n611));
  INV_X1    g425(.A(new_n383), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n436), .A2(new_n308), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n384), .B2(new_n436), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n325), .A2(new_n612), .A3(new_n454), .A4(new_n616), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n503), .A2(new_n560), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n617), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n562), .B1(new_n594), .B2(new_n596), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n591), .A2(new_n592), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n589), .B2(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n591), .A2(new_n592), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n627), .A2(G478), .A3(new_n308), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n553), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  AOI21_X1  g450(.A(new_n553), .B1(new_n597), .B2(new_n599), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n359), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n381), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n379), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n482), .A2(new_n496), .A3(new_n494), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n496), .B1(new_n482), .B2(new_n494), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n644), .B(new_n501), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n454), .A2(new_n325), .A3(new_n616), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n601), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT37), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G110), .ZN(G12));
  AOI21_X1  g466(.A(new_n647), .B1(new_n438), .B2(new_n450), .ZN(new_n653));
  INV_X1    g467(.A(new_n553), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n557), .B1(G900), .B2(new_n559), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n654), .A2(new_n600), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n325), .A2(new_n454), .A3(new_n653), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT98), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n201), .ZN(G30));
  NAND2_X1  g473(.A1(new_n325), .A2(new_n454), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n655), .B(KEYINPUT39), .Z(new_n661));
  OR3_X1    g475(.A1(new_n660), .A2(KEYINPUT40), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n411), .A2(new_n429), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n402), .A2(new_n439), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n308), .B1(new_n664), .B2(new_n416), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n438), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n644), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT40), .B1(new_n660), .B2(new_n661), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n645), .A2(new_n646), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n553), .A2(new_n501), .A3(new_n600), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n662), .A2(new_n668), .A3(new_n669), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  NAND3_X1  g489(.A1(new_n553), .A2(new_n631), .A3(new_n655), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n325), .A2(new_n454), .A3(new_n653), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  INV_X1    g493(.A(G469), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n302), .B2(new_n306), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n311), .B(new_n454), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n502), .A2(new_n561), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n451), .A3(new_n633), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n683), .A2(KEYINPUT99), .A3(new_n451), .A4(new_n633), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT41), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G113), .ZN(G15));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n451), .A3(new_n637), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  INV_X1    g506(.A(new_n682), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n653), .A2(new_n601), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  INV_X1    g509(.A(new_n384), .ZN(new_n696));
  INV_X1    g510(.A(new_n423), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n417), .B1(new_n429), .B2(new_n444), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n444), .A2(new_n429), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT100), .B1(new_n701), .B2(new_n417), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n696), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n383), .A3(new_n615), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n553), .A3(new_n600), .A4(new_n683), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND2_X1  g520(.A1(new_n700), .A2(new_n702), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n615), .B1(new_n707), .B2(new_n384), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n502), .A2(new_n682), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n644), .A3(new_n677), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(new_n501), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n605), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n498), .A2(new_n499), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n315), .A2(KEYINPUT101), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n297), .B1(new_n257), .B2(new_n255), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n312), .A4(new_n313), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(G469), .A3(new_n317), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(G469), .A2(G902), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n311), .A3(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n719), .A2(new_n311), .A3(KEYINPUT102), .A4(new_n720), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n714), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT103), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  MUX2_X1   g541(.A(new_n437), .B(new_n438), .S(new_n727), .Z(new_n728));
  AOI21_X1  g542(.A(new_n383), .B1(new_n728), .B2(new_n450), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n677), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n724), .ZN(new_n731));
  INV_X1    g545(.A(new_n714), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT103), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n734), .B(new_n714), .C1(new_n723), .C2(new_n724), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n451), .B(new_n677), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  OAI211_X1 g554(.A(new_n451), .B(new_n656), .C1(new_n733), .C2(new_n735), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  NOR2_X1   g556(.A1(new_n500), .A2(new_n712), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n631), .A2(new_n547), .A3(new_n551), .A4(new_n552), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT43), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n616), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n644), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT43), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n745), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n751), .B2(KEYINPUT105), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT106), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n752), .A3(new_n756), .A4(KEYINPUT44), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n744), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n754), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n320), .A2(new_n321), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(KEYINPUT45), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n317), .A4(new_n718), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(G469), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n720), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(KEYINPUT46), .B(new_n720), .C1(new_n764), .C2(new_n766), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n311), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n454), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n661), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n758), .A2(KEYINPUT107), .A3(new_n759), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n762), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n771), .A2(new_n778), .A3(new_n454), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n778), .B1(new_n771), .B2(new_n454), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n781), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT47), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n438), .A2(new_n450), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n612), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n744), .A2(new_n676), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n782), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  AND2_X1   g603(.A1(new_n667), .A2(new_n612), .ZN(new_n790));
  INV_X1    g604(.A(new_n311), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n681), .A2(new_n680), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT49), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n745), .A2(new_n712), .A3(new_n605), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(new_n794), .A3(new_n671), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n746), .A2(new_n557), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n704), .A3(new_n671), .A4(new_n693), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(new_n501), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT50), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n800), .B(KEYINPUT50), .C1(new_n798), .C2(new_n501), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n744), .A2(new_n682), .ZN(new_n805));
  INV_X1    g619(.A(new_n557), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n790), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n631), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n654), .A3(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n797), .A2(new_n704), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n743), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT113), .Z(new_n814));
  AOI22_X1  g628(.A1(new_n782), .A2(new_n784), .B1(new_n605), .B2(new_n793), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n804), .B(new_n811), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n797), .A2(new_n805), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n708), .A2(new_n644), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n816), .B2(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n809), .A2(new_n633), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n812), .A2(new_n503), .A3(new_n693), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n554), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n729), .A2(new_n797), .A3(new_n805), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n827), .A2(new_n828), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n822), .A2(new_n824), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n830), .A2(new_n831), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n657), .A2(new_n678), .A3(new_n710), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n500), .A2(new_n501), .A3(new_n553), .A4(new_n600), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n723), .B2(new_n724), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n379), .A2(new_n454), .A3(new_n643), .A4(new_n655), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n438), .B2(new_n666), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n841), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n672), .A2(new_n670), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n845), .A2(new_n731), .A3(new_n847), .A4(new_n841), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n839), .A2(new_n840), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n657), .A2(new_n678), .A3(new_n710), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n845), .A2(new_n731), .A3(new_n847), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT52), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n856), .A3(KEYINPUT111), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT109), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n597), .A2(new_n861), .A3(new_n599), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n597), .B2(new_n599), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n547), .A2(new_n551), .A3(new_n552), .A4(new_n655), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n644), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n714), .B1(new_n868), .B2(KEYINPUT110), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n867), .A2(new_n785), .A3(new_n869), .A4(new_n325), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n703), .A2(new_n749), .A3(new_n676), .A4(new_n615), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n733), .B2(new_n735), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n741), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n739), .A2(new_n851), .A3(new_n856), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n864), .A2(new_n654), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n632), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n617), .A2(new_n620), .A3(new_n622), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n691), .A2(new_n694), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n686), .B2(new_n687), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n649), .A2(new_n601), .B1(new_n455), .B2(new_n602), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n880), .A4(new_n705), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n859), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n739), .A2(new_n851), .A3(new_n856), .A4(new_n873), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n858), .B(new_n857), .C1(new_n884), .C2(new_n881), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n838), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n851), .A2(new_n856), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n741), .A2(new_n870), .A3(new_n872), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n738), .B2(new_n730), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n882), .A2(new_n887), .A3(new_n858), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT53), .B1(new_n884), .B2(new_n881), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT54), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR4_X1   g706(.A1(new_n836), .A2(new_n837), .A3(new_n886), .A4(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n796), .B1(new_n893), .B2(new_n894), .ZN(G75));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n891), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n308), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(G210), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n476), .B(new_n481), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n901), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n360), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  NOR4_X1   g719(.A1(new_n896), .A2(new_n308), .A3(new_n764), .A4(new_n766), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n720), .B(KEYINPUT57), .Z(new_n907));
  NAND3_X1  g721(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT54), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n892), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n910), .B2(new_n307), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT117), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  INV_X1    g727(.A(new_n904), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n896), .A2(new_n838), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n908), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n916), .A2(new_n907), .B1(new_n306), .B2(new_n302), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n913), .B(new_n914), .C1(new_n917), .C2(new_n906), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n543), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n904), .ZN(G60));
  AND2_X1   g738(.A1(new_n627), .A2(new_n629), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT118), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT59), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n916), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n886), .B2(new_n892), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n931), .A2(new_n932), .A3(new_n926), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n931), .B2(new_n926), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n914), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(G63));
  INV_X1    g750(.A(new_n896), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT120), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n380), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n642), .A3(new_n940), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n914), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G66));
  AOI21_X1  g760(.A(new_n360), .B1(new_n558), .B2(G224), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n881), .B2(new_n360), .ZN(new_n948));
  INV_X1    g762(.A(G898), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n476), .B1(new_n949), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT121), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n948), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(G900), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n299), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT124), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n729), .A2(new_n847), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n758), .A2(KEYINPUT107), .A3(new_n759), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT107), .B1(new_n758), .B2(new_n759), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n773), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n788), .A2(new_n739), .A3(new_n839), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n360), .A3(new_n741), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n410), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(G900), .A2(G953), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n788), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n958), .A2(new_n959), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n773), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n674), .B2(new_n839), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(KEYINPUT123), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n660), .A2(new_n661), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n451), .A3(new_n743), .A4(new_n876), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n674), .A2(new_n972), .A3(new_n839), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT122), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n971), .A2(new_n976), .A3(new_n978), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n966), .B1(new_n982), .B2(new_n360), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n956), .B1(new_n968), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n775), .A2(new_n788), .A3(new_n978), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n974), .A2(new_n975), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n986), .A3(new_n980), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n965), .B1(new_n987), .B2(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n955), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n984), .A2(new_n990), .ZN(G72));
  INV_X1    g805(.A(new_n411), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n961), .A2(new_n741), .A3(new_n882), .A4(new_n962), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT125), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT63), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n992), .B(new_n416), .C1(new_n993), .C2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n663), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n775), .A2(new_n788), .A3(new_n978), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(new_n882), .A3(new_n976), .A4(new_n981), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n1001), .B2(new_n997), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n883), .A2(new_n885), .ZN(new_n1003));
  INV_X1    g817(.A(new_n434), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1003), .B(new_n997), .C1(new_n1004), .C2(new_n447), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n914), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n998), .A2(new_n1002), .A3(new_n1006), .ZN(G57));
endmodule


