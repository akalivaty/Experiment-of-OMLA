//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G77), .A2(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n209), .B(new_n213), .C1(G50), .C2(G226), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G97), .A2(G257), .ZN(new_n216));
  XOR2_X1   g0016(.A(KEYINPUT65), .B(G238), .Z(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n206), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n224), .B(new_n227), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n204), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n228), .B1(new_n230), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n208), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G179), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  OAI211_X1 g0053(.A(G1), .B(G13), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT69), .B1(new_n254), .B2(new_n255), .ZN(new_n259));
  OAI21_X1  g0059(.A(G238), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n252), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n212), .A2(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G226), .B2(G1698), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n261), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n255), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n260), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT72), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n260), .A2(new_n278), .A3(new_n271), .A4(new_n274), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n251), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n276), .A2(new_n279), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G169), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  AOI211_X1 g0088(.A(new_n288), .B(new_n284), .C1(new_n276), .C2(new_n279), .ZN(new_n289));
  OR3_X1    g0089(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n229), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n204), .A2(G1), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT12), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n218), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n204), .A2(G33), .A3(G77), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G50), .ZN(new_n304));
  OAI221_X1 g0104(.A(new_n301), .B1(new_n204), .B2(G68), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n295), .ZN(new_n306));
  XOR2_X1   g0106(.A(new_n306), .B(KEYINPUT11), .Z(new_n307));
  INV_X1    g0107(.A(new_n291), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(KEYINPUT12), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n300), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n293), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n311), .A2(new_n298), .A3(G68), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n291), .A2(G50), .ZN(new_n316));
  NOR4_X1   g0116(.A1(new_n308), .A2(new_n295), .A3(new_n304), .A4(new_n296), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(G20), .A3(new_n252), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  NOR3_X1   g0120(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n320), .A2(new_n303), .B1(new_n321), .B2(new_n204), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n295), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT70), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(new_n295), .C1(new_n319), .C2(new_n322), .ZN(new_n326));
  AOI211_X1 g0126(.A(new_n316), .B(new_n317), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n256), .B(new_n257), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G226), .ZN(new_n329));
  INV_X1    g0129(.A(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G222), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G223), .A2(G1698), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n265), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n333), .B(new_n270), .C1(G77), .C2(new_n265), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n329), .A2(new_n274), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G179), .ZN(new_n336));
  AOI211_X1 g0136(.A(new_n327), .B(new_n336), .C1(new_n288), .C2(new_n335), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(G200), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n329), .A2(G190), .A3(new_n274), .A4(new_n334), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n317), .B1(new_n324), .B2(new_n326), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(G50), .B2(new_n291), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT9), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n338), .B(new_n339), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n327), .A2(KEYINPUT9), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT10), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n339), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(KEYINPUT9), .B2(new_n327), .ZN(new_n347));
  INV_X1    g0147(.A(new_n344), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n337), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n314), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n280), .B2(new_n281), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n286), .A2(G200), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n273), .B1(new_n328), .B2(G244), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n217), .A2(new_n330), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n265), .B1(new_n212), .B2(G1698), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n359), .A2(new_n360), .B1(G107), .B2(new_n265), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n254), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT15), .B(G87), .Z(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n204), .A3(G33), .ZN(new_n365));
  INV_X1    g0165(.A(G77), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n365), .B1(new_n204), .B2(new_n366), .C1(new_n303), .C2(new_n318), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n295), .B1(new_n297), .B2(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n293), .A2(new_n366), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n363), .B(new_n371), .C1(new_n353), .C2(new_n362), .ZN(new_n372));
  AND4_X1   g0172(.A1(new_n315), .A2(new_n351), .A3(new_n357), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n264), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(G226), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n265), .A2(new_n378), .A3(G226), .A4(G1698), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n265), .A2(G223), .A3(new_n330), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n273), .B1(new_n382), .B2(new_n270), .ZN(new_n383));
  OR2_X1    g0183(.A1(KEYINPUT77), .A2(G190), .ZN(new_n384));
  NAND2_X1  g0184(.A1(KEYINPUT77), .A2(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n256), .A2(new_n212), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AOI211_X1 g0189(.A(new_n273), .B(new_n387), .C1(new_n382), .C2(new_n270), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(G200), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT75), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n263), .A2(new_n204), .A3(new_n264), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n264), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT74), .A3(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G68), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n211), .A2(new_n218), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n302), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n218), .B1(new_n395), .B2(new_n396), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n295), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n392), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n318), .A2(new_n296), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n308), .A2(new_n295), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n412), .A2(new_n413), .B1(new_n308), .B2(new_n318), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(KEYINPUT75), .A3(new_n295), .A4(new_n409), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n391), .A2(new_n411), .A3(new_n414), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n411), .A2(new_n416), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n420), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n391), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n390), .A2(G179), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n288), .B2(new_n390), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n422), .A2(KEYINPUT18), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT18), .B1(new_n422), .B2(new_n424), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n419), .B(new_n421), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n362), .A2(G179), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n362), .A2(new_n288), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n370), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT78), .B1(new_n373), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n315), .A2(new_n351), .A3(new_n357), .A4(new_n372), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n425), .A2(new_n426), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(new_n419), .A3(new_n421), .A4(new_n430), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n265), .A2(G244), .A3(new_n330), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT4), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n265), .A2(new_n444), .A3(G244), .A4(new_n330), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n270), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(new_n272), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n254), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G257), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n451), .A2(new_n251), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n295), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT6), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(G97), .A2(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n470), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n395), .A2(new_n396), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n462), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n413), .B1(G1), .B2(new_n252), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n464), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n291), .A2(G97), .ZN(new_n477));
  OR3_X1    g0277(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n457), .ZN(new_n479));
  INV_X1    g0279(.A(new_n460), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n479), .B(new_n480), .C1(new_n450), .C2(new_n270), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n461), .B(new_n478), .C1(new_n481), .C2(G169), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n453), .A2(G250), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n270), .B(new_n483), .C1(new_n272), .C2(new_n453), .ZN(new_n484));
  OR2_X1    g0284(.A1(G238), .A2(G1698), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n265), .B(new_n485), .C1(G244), .C2(new_n330), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G116), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n254), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G190), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n265), .A2(new_n204), .A3(G68), .ZN(new_n491));
  INV_X1    g0291(.A(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n467), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n261), .A2(new_n204), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(KEYINPUT19), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n261), .A2(G20), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n491), .B(new_n495), .C1(KEYINPUT19), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n295), .ZN(new_n498));
  INV_X1    g0298(.A(new_n364), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n293), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n475), .A2(new_n492), .ZN(new_n502));
  OAI21_X1  g0302(.A(G200), .B1(new_n484), .B2(new_n488), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n490), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n498), .B(new_n500), .C1(new_n499), .C2(new_n475), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n489), .A2(new_n251), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n288), .B1(new_n484), .B2(new_n488), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n451), .A2(G190), .A3(new_n457), .A4(new_n460), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n512));
  INV_X1    g0312(.A(G200), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n511), .B(new_n512), .C1(new_n481), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n265), .A2(G250), .A3(new_n330), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT84), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT84), .A4(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n270), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n459), .A2(G264), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n457), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n413), .B(G107), .C1(G1), .C2(new_n252), .ZN(new_n526));
  INV_X1    g0326(.A(G13), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G1), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n204), .A2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT82), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT25), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n531), .A2(KEYINPUT25), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(KEYINPUT25), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n533), .A2(new_n528), .A3(new_n534), .A4(new_n529), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n526), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n526), .A2(KEYINPUT83), .A3(new_n532), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n265), .A2(new_n204), .A3(G87), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n529), .A2(KEYINPUT23), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n541), .A2(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n265), .A2(new_n547), .A3(new_n204), .A4(G87), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT24), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n546), .A2(KEYINPUT24), .A3(new_n548), .A4(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n295), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n522), .A2(G190), .A3(new_n457), .A4(new_n523), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n525), .A2(new_n540), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  AND4_X1   g0356(.A1(new_n482), .A2(new_n510), .A3(new_n514), .A4(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n207), .B1(new_n203), .B2(G33), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n311), .A2(new_n462), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n293), .A2(new_n207), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n447), .B(new_n204), .C1(G33), .C2(new_n464), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n561), .B(new_n295), .C1(new_n204), .C2(G116), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n559), .B(new_n560), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n457), .B1(new_n208), .B2(new_n458), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n265), .A2(G264), .A3(G1698), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n265), .A2(G257), .A3(new_n330), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT80), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n265), .A2(new_n571), .A3(G264), .A4(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n266), .A2(G303), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n569), .A2(new_n570), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n567), .B1(new_n574), .B2(new_n270), .ZN(new_n575));
  INV_X1    g0375(.A(new_n386), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n566), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n513), .B2(new_n575), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n554), .A2(new_n540), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n524), .A2(new_n288), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n522), .A2(new_n251), .A3(new_n457), .A4(new_n523), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(G179), .A3(new_n566), .ZN(new_n583));
  INV_X1    g0383(.A(new_n575), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(G169), .A3(new_n566), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n584), .A2(KEYINPUT21), .A3(G169), .A4(new_n566), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n582), .A2(new_n583), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n557), .A2(new_n578), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n439), .A2(new_n591), .ZN(G372));
  AOI22_X1  g0392(.A1(new_n314), .A2(new_n290), .B1(new_n357), .B2(new_n431), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n421), .A2(new_n419), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n435), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n345), .A2(new_n350), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n337), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n587), .A2(new_n588), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT85), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n583), .A4(new_n582), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n557), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n508), .ZN(new_n603));
  INV_X1    g0403(.A(new_n482), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(KEYINPUT26), .A3(new_n510), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT26), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n482), .B2(new_n509), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n603), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n597), .B1(new_n439), .B2(new_n609), .ZN(G369));
  NAND3_X1  g0410(.A1(new_n587), .A2(new_n583), .A3(new_n588), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n528), .A2(new_n204), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(G213), .ZN(new_n615));
  INV_X1    g0415(.A(G343), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n566), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n578), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G330), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n579), .A2(new_n617), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n556), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n582), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n582), .B2(new_n617), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n617), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n582), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT86), .ZN(G399));
  INV_X1    g0437(.A(new_n225), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(G41), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n493), .A2(G116), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G1), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n232), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n640), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT28), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n557), .A2(new_n589), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n617), .B1(new_n608), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT29), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT29), .B(new_n617), .C1(new_n602), .C2(new_n608), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n574), .A2(new_n270), .ZN(new_n652));
  INV_X1    g0452(.A(new_n567), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(G179), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n522), .A2(new_n523), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(new_n481), .A3(KEYINPUT30), .A4(new_n489), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT30), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n451), .A2(new_n457), .A3(new_n460), .A4(new_n489), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n575), .A2(G179), .A3(new_n523), .A4(new_n522), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n451), .A2(new_n457), .A3(new_n460), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(new_n251), .A3(new_n584), .A4(new_n524), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n657), .B(new_n661), .C1(new_n489), .C2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n664), .A2(KEYINPUT31), .A3(new_n617), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT31), .B1(new_n664), .B2(new_n617), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT87), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n617), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT31), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT87), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n664), .A2(KEYINPUT31), .A3(new_n617), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n557), .A2(new_n578), .A3(new_n590), .A4(new_n631), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n651), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n645), .B1(new_n678), .B2(G1), .ZN(G364));
  AOI21_X1  g0479(.A(new_n229), .B1(G20), .B2(new_n288), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n204), .A2(new_n251), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G200), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G190), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(KEYINPUT33), .A2(G317), .ZN(new_n685));
  NOR2_X1   g0485(.A1(KEYINPUT33), .A2(G317), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n251), .A2(G200), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n689), .A2(new_n204), .A3(new_n353), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n265), .B1(new_n690), .B2(G303), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT96), .Z(new_n692));
  INV_X1    g0492(.A(G283), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(G20), .B2(new_n353), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n204), .A2(KEYINPUT92), .A3(G190), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n689), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n697), .A2(G179), .A3(G200), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G329), .ZN(new_n704));
  OAI221_X1 g0504(.A(new_n692), .B1(new_n693), .B2(new_n699), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n681), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n707), .A2(new_n513), .A3(new_n576), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n688), .B(new_n705), .C1(G322), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G294), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G179), .A2(G200), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n204), .B1(new_n712), .B2(G190), .ZN(new_n713));
  INV_X1    g0513(.A(G311), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n353), .A3(new_n513), .ZN(new_n715));
  OAI221_X1 g0515(.A(new_n710), .B1(new_n711), .B2(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n682), .A2(new_n386), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(G326), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT93), .B(G159), .Z(new_n720));
  NAND2_X1  g0520(.A1(new_n700), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT94), .Z(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT32), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n709), .A2(G58), .B1(G107), .B2(new_n698), .ZN(new_n724));
  INV_X1    g0524(.A(new_n715), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G77), .ZN(new_n726));
  INV_X1    g0526(.A(new_n713), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G97), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n723), .A2(new_n724), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n690), .A2(G87), .ZN(new_n730));
  INV_X1    g0530(.A(new_n717), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(new_n304), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n722), .A2(KEYINPUT32), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n265), .B1(new_n684), .B2(new_n218), .ZN(new_n734));
  NOR4_X1   g0534(.A1(new_n729), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT95), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n680), .B1(new_n719), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n527), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n640), .A2(G1), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n621), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n638), .A2(new_n207), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n249), .A2(new_n452), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n638), .A2(new_n265), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n643), .B2(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n225), .A2(new_n265), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT89), .Z(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(G355), .B(KEYINPUT90), .Z(new_n753));
  OAI221_X1 g0553(.A(new_n746), .B1(new_n747), .B2(new_n749), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n744), .A2(new_n680), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n737), .A2(new_n741), .A3(new_n745), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n621), .A2(new_n622), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n624), .A2(new_n740), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(G396));
  NAND2_X1  g0560(.A1(new_n698), .A2(G87), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n703), .B2(new_n714), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT98), .Z(new_n763));
  OAI21_X1  g0563(.A(new_n266), .B1(new_n715), .B2(new_n207), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n728), .B1(new_n731), .B2(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n683), .A2(G283), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n690), .A2(G107), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n709), .A2(G294), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n709), .A2(G143), .B1(G150), .B2(new_n683), .ZN(new_n772));
  INV_X1    g0572(.A(G137), .ZN(new_n773));
  INV_X1    g0573(.A(new_n720), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n772), .B1(new_n773), .B2(new_n731), .C1(new_n715), .C2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT34), .ZN(new_n777));
  INV_X1    g0577(.A(new_n703), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n266), .B1(new_n778), .B2(G132), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n698), .A2(G68), .B1(G58), .B2(new_n727), .ZN(new_n780));
  INV_X1    g0580(.A(new_n690), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n779), .B(new_n780), .C1(new_n304), .C2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n771), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n372), .B1(new_n371), .B2(new_n631), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n430), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n431), .A2(new_n631), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n783), .A2(new_n680), .B1(new_n742), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n680), .A2(new_n742), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n741), .C1(G77), .C2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT100), .Z(new_n792));
  NOR2_X1   g0592(.A1(new_n609), .A2(new_n617), .ZN(new_n793));
  INV_X1    g0593(.A(new_n787), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n787), .B1(new_n609), .B2(new_n617), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n795), .A2(G330), .A3(new_n675), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n740), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(KEYINPUT101), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n676), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT101), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n797), .A2(new_n802), .A3(new_n740), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(new_n804), .ZN(G384));
  NAND3_X1  g0605(.A1(new_n674), .A2(new_n670), .A3(new_n672), .ZN(new_n806));
  INV_X1    g0606(.A(new_n356), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n314), .A2(new_n807), .A3(new_n354), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n314), .B(new_n617), .C1(new_n290), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n314), .A2(new_n617), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n357), .B(new_n810), .C1(new_n811), .C2(new_n352), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n806), .A2(new_n813), .A3(new_n794), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT103), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n615), .B(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n422), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n427), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n815), .B1(new_n427), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n422), .A2(new_n424), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n817), .A3(new_n417), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT37), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n817), .A3(new_n825), .A4(new_n417), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT38), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n415), .A2(new_n295), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT16), .B1(new_n399), .B2(new_n405), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n414), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n615), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n427), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n831), .B1(new_n424), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n417), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n826), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n427), .A2(new_n833), .B1(new_n837), .B2(new_n826), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(KEYINPUT104), .A3(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT40), .B(new_n814), .C1(new_n828), .C2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n839), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n842), .A2(KEYINPUT38), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n814), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT40), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(new_n850), .A3(G330), .ZN(new_n851));
  OAI211_X1 g0651(.A(G330), .B(new_n806), .C1(new_n433), .C2(new_n438), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT106), .Z(new_n854));
  OAI21_X1  g0654(.A(new_n806), .B1(new_n433), .B2(new_n438), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n845), .A2(new_n850), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n433), .A2(new_n438), .B1(new_n649), .B2(new_n650), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n597), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n857), .B(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n425), .A2(new_n426), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n818), .B1(new_n861), .B2(new_n594), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT103), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n427), .A2(new_n815), .A3(new_n818), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n827), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT39), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n841), .A4(new_n843), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT105), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n846), .A2(new_n847), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  INV_X1    g0672(.A(new_n844), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n868), .A4(new_n867), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n315), .A2(new_n617), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n435), .A2(new_n816), .ZN(new_n879));
  INV_X1    g0679(.A(new_n786), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n793), .B2(new_n794), .ZN(new_n881));
  INV_X1    g0681(.A(new_n813), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n879), .B1(new_n883), .B2(new_n871), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n860), .B(new_n885), .Z(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n203), .B2(new_n738), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n207), .B1(new_n470), .B2(KEYINPUT35), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n888), .B(new_n230), .C1(KEYINPUT35), .C2(new_n470), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT36), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n643), .A2(new_n366), .A3(new_n400), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n218), .A2(G50), .ZN(new_n892));
  OAI211_X1 g0692(.A(G1), .B(new_n527), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n890), .A3(new_n893), .ZN(G367));
  NAND2_X1  g0694(.A1(new_n739), .A2(G1), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n604), .A2(new_n617), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n482), .B(new_n514), .C1(new_n512), .C2(new_n631), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n635), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT45), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n635), .A2(KEYINPUT44), .A3(new_n898), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT44), .B1(new_n635), .B2(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n900), .A2(new_n903), .A3(new_n629), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n629), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n628), .A2(new_n632), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n908), .A2(KEYINPUT108), .A3(new_n633), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT108), .B1(new_n908), .B2(new_n633), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n623), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n910), .A2(new_n623), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n678), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n639), .B(KEYINPUT41), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n895), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n629), .A2(new_n898), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n631), .B1(new_n501), .B2(new_n502), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n603), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n509), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT107), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n918), .B(new_n923), .Z(new_n924));
  NAND2_X1  g0724(.A1(new_n633), .A2(new_n898), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT42), .Z(new_n926));
  OAI21_X1  g0726(.A(new_n482), .B1(new_n897), .B2(new_n582), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n631), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n926), .A2(new_n928), .B1(KEYINPUT43), .B2(new_n921), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n924), .B(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n921), .A2(G20), .A3(new_n743), .ZN(new_n931));
  INV_X1    g0731(.A(new_n748), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n755), .B1(new_n225), .B2(new_n499), .C1(new_n236), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n700), .A2(G317), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n465), .B2(new_n713), .C1(new_n714), .C2(new_n731), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT46), .B1(new_n690), .B2(G116), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(G294), .B2(new_n683), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n265), .B1(new_n698), .B2(G97), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n690), .A2(KEYINPUT46), .A3(G116), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n715), .A2(new_n693), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n708), .A2(new_n765), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n935), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n266), .B1(new_n727), .B2(G68), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n699), .B2(new_n366), .C1(new_n304), .C2(new_n715), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n709), .A2(G150), .B1(G137), .B2(new_n700), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n684), .B2(new_n774), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n945), .B(new_n947), .C1(G143), .C2(new_n717), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n690), .A2(G58), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g0752(.A(new_n680), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n741), .B(new_n933), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n917), .A2(new_n930), .B1(new_n931), .B2(new_n954), .ZN(G387));
  OR2_X1    g0755(.A1(new_n678), .A2(new_n913), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n678), .A2(new_n913), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n639), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n748), .B1(new_n241), .B2(new_n452), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n752), .B2(new_n641), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n318), .A2(G50), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT50), .ZN(new_n962));
  AOI21_X1  g0762(.A(G45), .B1(G68), .B2(G77), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n641), .A3(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n960), .A2(new_n964), .B1(new_n465), .B2(new_n638), .ZN(new_n965));
  INV_X1    g0765(.A(new_n755), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n741), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n709), .A2(G317), .B1(G311), .B2(new_n683), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n717), .A2(G322), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n765), .C2(new_n715), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n693), .B2(new_n713), .C1(new_n711), .C2(new_n781), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT49), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n265), .B1(new_n700), .B2(G326), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n207), .C2(new_n699), .ZN(new_n975));
  INV_X1    g0775(.A(G159), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n731), .A2(new_n976), .B1(new_n684), .B2(new_n318), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n265), .B1(new_n715), .B2(new_n218), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(new_n364), .C2(new_n727), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n700), .A2(G150), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n366), .B2(new_n781), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n709), .A2(G50), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n981), .A2(KEYINPUT110), .B1(G97), .B2(new_n698), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n953), .B1(new_n975), .B2(new_n985), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n967), .B(new_n986), .C1(new_n628), .C2(new_n744), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n913), .B2(new_n895), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n958), .A2(new_n988), .ZN(G393));
  AOI21_X1  g0789(.A(new_n640), .B1(new_n906), .B2(new_n957), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n906), .B2(new_n957), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n904), .A2(new_n895), .A3(new_n905), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n709), .A2(G311), .B1(G317), .B2(new_n717), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT52), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n698), .A2(G107), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n690), .A2(G283), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n700), .A2(G322), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n684), .A2(new_n765), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n713), .A2(new_n207), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n266), .B1(new_n715), .B2(new_n711), .ZN(new_n1001));
  NOR4_X1   g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n708), .A2(new_n976), .B1(new_n320), .B2(new_n731), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT51), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n727), .A2(G77), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n700), .A2(G143), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n761), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n684), .A2(new_n304), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n781), .A2(new_n218), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n265), .B1(new_n715), .B2(new_n318), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n680), .B1(new_n1002), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n896), .A2(new_n897), .A3(new_n744), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n966), .B1(new_n748), .B2(new_n245), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n464), .B2(new_n225), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n741), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n991), .A2(new_n992), .A3(new_n1016), .ZN(G390));
  XOR2_X1   g0817(.A(KEYINPUT54), .B(G143), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n725), .A2(new_n1018), .B1(G137), .B2(new_n683), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT112), .Z(new_n1020));
  NAND2_X1  g0820(.A1(new_n690), .A2(G150), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT53), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n778), .A2(G125), .ZN(new_n1023));
  INV_X1    g0823(.A(G132), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n265), .B1(new_n699), .B2(new_n304), .C1(new_n708), .C2(new_n1024), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(G128), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n731), .C1(new_n976), .C2(new_n713), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n730), .B1(new_n465), .B2(new_n684), .C1(new_n715), .C2(new_n464), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G68), .B2(new_n698), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n266), .B(new_n1005), .C1(new_n731), .C2(new_n693), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n709), .B2(G116), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(new_n711), .C2(new_n703), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n680), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n876), .B2(new_n743), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n789), .A2(new_n318), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1036), .A2(new_n740), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT113), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n877), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n881), .B2(new_n882), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n870), .A2(new_n1042), .A3(new_n875), .A4(new_n872), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n880), .B1(new_n647), .B2(new_n785), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1041), .B1(new_n882), .B2(new_n1044), .C1(new_n828), .C2(new_n844), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n675), .A2(G330), .A3(new_n794), .A4(new_n813), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n806), .A2(new_n813), .A3(G330), .A4(new_n794), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n895), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n852), .A2(new_n858), .A3(new_n597), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n806), .A2(G330), .A3(new_n794), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n882), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT111), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1059), .A3(new_n882), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1058), .A2(new_n1044), .A3(new_n1046), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n675), .A2(G330), .A3(new_n794), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1051), .B1(new_n1063), .B2(new_n882), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(new_n881), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1055), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1052), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1069), .A2(new_n1048), .A3(new_n1066), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1070), .A3(new_n639), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1040), .A2(new_n1053), .A3(new_n1071), .ZN(G378));
  NOR2_X1   g0872(.A1(new_n790), .A2(G50), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n698), .A2(G58), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n253), .C1(new_n207), .C2(new_n731), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n727), .A2(G68), .B1(new_n690), .B2(G77), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n265), .B1(new_n683), .B2(G97), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n708), .C2(new_n465), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1075), .B(new_n1078), .C1(new_n364), .C2(new_n725), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n693), .B2(new_n703), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT58), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n304), .B1(new_n374), .B2(G41), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n709), .A2(G128), .B1(new_n690), .B2(new_n1018), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n725), .A2(G137), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n717), .A2(G125), .B1(G150), .B2(new_n727), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G132), .B2(new_n683), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT59), .ZN(new_n1088));
  AOI21_X1  g0888(.A(G41), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n698), .A2(new_n720), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT114), .B(G124), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n700), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n252), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1081), .B(new_n1082), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n740), .B(new_n1073), .C1(new_n1095), .C2(new_n680), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n351), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n351), .A2(new_n1097), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n327), .A2(new_n615), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1096), .B1(new_n1109), .B2(new_n743), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1109), .A2(new_n845), .A3(G330), .A4(new_n850), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n851), .A2(new_n1113), .ZN(new_n1114));
  AND4_X1   g0914(.A1(new_n878), .A2(new_n884), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n878), .A2(new_n884), .B1(new_n1114), .B2(new_n1112), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT116), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n885), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1111), .B1(new_n1122), .B2(new_n895), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1068), .A2(new_n1055), .ZN(new_n1124));
  AOI21_X1  g0924(.A(KEYINPUT57), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n878), .A2(new_n884), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n639), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1123), .B1(new_n1125), .B2(new_n1130), .ZN(G375));
  NAND2_X1  g0931(.A1(new_n1063), .A2(new_n882), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1050), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n881), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n1061), .B1(G1), .B2(new_n739), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n731), .A2(new_n711), .B1(new_n499), .B2(new_n713), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n265), .B1(new_n698), .B2(G77), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT118), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n693), .B2(new_n708), .C1(new_n765), .C2(new_n703), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(G107), .C2(new_n725), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n464), .B2(new_n781), .C1(new_n207), .C2(new_n684), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT119), .Z(new_n1143));
  AOI22_X1  g0943(.A1(new_n778), .A2(G128), .B1(G137), .B2(new_n709), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n717), .A2(G132), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1074), .B1(new_n304), .B2(new_n713), .C1(new_n715), .C2(new_n320), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G159), .B2(new_n690), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n265), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n683), .B2(new_n1018), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n680), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n882), .A2(new_n742), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n740), .B1(new_n218), .B2(new_n789), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT117), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT120), .B1(new_n1136), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n895), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT120), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1054), .B(new_n1061), .C1(new_n881), .C2(new_n1064), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1066), .A2(new_n916), .A3(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(G381));
  NOR2_X1   g0964(.A1(G387), .A2(G384), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n1163), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT121), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n640), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1117), .A2(new_n1121), .B1(new_n1055), .B2(new_n1068), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(KEYINPUT57), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1040), .A2(new_n1053), .A3(new_n1071), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1123), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1165), .A2(new_n1166), .A3(KEYINPUT121), .A4(new_n1163), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1169), .A2(new_n1175), .A3(new_n1176), .ZN(G407));
  INV_X1    g0977(.A(G213), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(G343), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR3_X1    g0980(.A1(new_n1174), .A2(KEYINPUT122), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT122), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(G407), .A2(new_n1181), .A3(G213), .A4(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT123), .Z(G409));
  INV_X1    g0984(.A(KEYINPUT126), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1161), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1135), .A2(KEYINPUT60), .A3(new_n1061), .A4(new_n1054), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1187), .A2(new_n639), .A3(new_n1066), .A4(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1136), .A2(KEYINPUT120), .A3(new_n1155), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1158), .B1(new_n1157), .B2(new_n1154), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1189), .B(G384), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G384), .B1(new_n1160), .B2(new_n1189), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT124), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1179), .A2(G2897), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1197));
  INV_X1    g0997(.A(G384), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n1192), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1196), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1203), .A2(new_n1200), .A3(G2897), .A4(new_n1179), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1179), .B1(G375), .B2(G378), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1120), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1124), .B(new_n916), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n895), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1110), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(G378), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1205), .B1(new_n1206), .B2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1185), .B1(new_n1214), .B2(KEYINPUT61), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT61), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1173), .B1(new_n1172), .B2(new_n1123), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1217), .A2(new_n1212), .A3(new_n1179), .ZN(new_n1218));
  OAI211_X1 g1018(.A(KEYINPUT126), .B(new_n1216), .C1(new_n1218), .C2(new_n1205), .ZN(new_n1219));
  AND2_X1   g1019(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1218), .A2(new_n1203), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1203), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1215), .A2(new_n1219), .A3(new_n1223), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(G387), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(G387), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1228), .B2(G387), .ZN(new_n1234));
  XOR2_X1   g1034(.A(G393), .B(G396), .Z(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1232), .B(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1227), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT63), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1224), .A2(new_n1239), .A3(new_n1225), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(new_n1237), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1214), .A2(new_n1239), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n1216), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1238), .A2(new_n1243), .ZN(G405));
  OR2_X1    g1044(.A1(new_n1175), .A2(new_n1217), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1225), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1237), .A2(new_n1245), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1203), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G402));
endmodule


