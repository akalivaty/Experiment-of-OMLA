//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G353));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n202), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n206), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n216), .B(new_n217), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n224), .B1(new_n223), .B2(new_n222), .C1(new_n209), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  NAND2_X1  g0029(.A1(new_n204), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n227), .A2(G13), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n236), .B(G250), .C1(G257), .C2(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT0), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n229), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(G361));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G250), .B(G257), .Z(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XOR2_X1   g0055(.A(KEYINPUT8), .B(G58), .Z(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .C1(new_n205), .C2(new_n233), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n232), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n219), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n265), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(G50), .C1(G1), .C2(new_n233), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT68), .B1(new_n277), .B2(new_n232), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(G1), .A4(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT66), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT66), .A2(G41), .ZN(new_n288));
  AOI21_X1  g0088(.A(G45), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT67), .B1(new_n289), .B2(G1), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n278), .B2(new_n281), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  INV_X1    g0093(.A(new_n288), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT66), .A2(G41), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n297), .A3(new_n267), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n290), .A2(new_n292), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT3), .B(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G222), .ZN(new_n302));
  INV_X1    g0102(.A(G223), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n300), .B(new_n302), .C1(new_n303), .C2(new_n301), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n277), .A2(new_n232), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n304), .B(new_n305), .C1(G77), .C2(new_n300), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n286), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G200), .ZN(new_n308));
  INV_X1    g0108(.A(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G190), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n275), .A2(new_n276), .A3(new_n308), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT10), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT69), .B(G179), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n273), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n303), .A2(new_n301), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n220), .A2(G1698), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n320), .A2(new_n321), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n257), .B2(new_n214), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n305), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n299), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n316), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n313), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n233), .B1(new_n204), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n300), .B2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n320), .A2(new_n323), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT7), .A3(new_n233), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n333), .B1(new_n338), .B2(G68), .ZN(new_n339));
  INV_X1    g0139(.A(G159), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n262), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT16), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n203), .B1(new_n335), .B2(new_n337), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NOR4_X1   g0145(.A1(new_n344), .A2(new_n345), .A3(new_n341), .A4(new_n333), .ZN(new_n346));
  INV_X1    g0146(.A(new_n265), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n343), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n256), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n267), .B2(G20), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n271), .B1(new_n269), .B2(new_n349), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n330), .B(new_n331), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT18), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT7), .B1(new_n336), .B2(new_n233), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n334), .B(G20), .C1(new_n320), .C2(new_n323), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n333), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n342), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n345), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n342), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n265), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n351), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT18), .A3(new_n330), .A4(new_n331), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n329), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n299), .A2(new_n327), .A3(new_n369), .A4(new_n328), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n363), .A2(new_n371), .A3(new_n351), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n363), .A2(new_n371), .A3(new_n351), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n299), .B1(new_n221), .B2(new_n284), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT70), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G238), .A2(G1698), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n300), .B(new_n382), .C1(new_n213), .C2(G1698), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n305), .C1(G107), .C2(new_n300), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G200), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n347), .B2(new_n268), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n269), .A2(new_n265), .A3(KEYINPUT71), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n267), .B2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n269), .A2(new_n206), .ZN(new_n393));
  XOR2_X1   g0193(.A(KEYINPUT15), .B(G87), .Z(new_n394));
  AOI22_X1  g0194(.A1(new_n261), .A2(new_n256), .B1(new_n394), .B2(new_n258), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n233), .B2(new_n206), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n265), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n381), .A2(G190), .A3(new_n384), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n386), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n366), .A2(new_n379), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n319), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(new_n385), .B2(new_n316), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n381), .A2(new_n314), .A3(new_n384), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n320), .A2(new_n323), .A3(G232), .A4(G1698), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n300), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n320), .A2(new_n323), .A3(G226), .A4(new_n301), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT73), .B1(new_n412), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(new_n305), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n285), .A2(G238), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n299), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT13), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n412), .A2(new_n415), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT73), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n415), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n305), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n420), .A4(new_n299), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n422), .A2(new_n423), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(KEYINPUT74), .B(KEYINPUT13), .C1(new_n419), .C2(new_n421), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(G169), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n422), .A2(G179), .A3(new_n430), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n431), .A2(new_n436), .A3(G169), .A4(new_n432), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n391), .A2(G68), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n258), .A2(G77), .B1(new_n261), .B2(G50), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n233), .B2(G68), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n265), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT11), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT12), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n269), .B(new_n203), .C1(KEYINPUT76), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(KEYINPUT76), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n439), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n407), .B1(new_n438), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n422), .A2(G190), .A3(new_n430), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n422), .A2(new_n430), .A3(KEYINPUT75), .A4(G190), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n448), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n431), .A2(G200), .A3(new_n432), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n403), .A2(new_n449), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n320), .A2(new_n323), .A3(G244), .A4(G1698), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n300), .A2(new_n462), .A3(G244), .A4(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G116), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n300), .A2(G238), .A3(new_n301), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n461), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n305), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n293), .A2(G1), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G250), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n278), .B2(new_n281), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n291), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n367), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n233), .A2(G33), .A3(G97), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT19), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n233), .B1(new_n414), .B2(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n214), .A2(new_n209), .A3(new_n210), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n320), .A2(new_n323), .A3(new_n233), .A4(G68), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n474), .A2(KEYINPUT82), .A3(new_n475), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n478), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n265), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n394), .A2(new_n268), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n267), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n268), .A2(new_n488), .A3(new_n232), .A4(new_n264), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n485), .B(new_n487), .C1(new_n214), .C2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n459), .B1(new_n473), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n466), .A2(new_n305), .B1(new_n470), .B2(new_n471), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n489), .A2(new_n214), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n486), .B(new_n494), .C1(new_n484), .C2(new_n265), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(KEYINPUT83), .C1(new_n492), .C2(new_n367), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n314), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n394), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n485), .B(new_n487), .C1(new_n501), .C2(new_n489), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n492), .A2(KEYINPUT81), .A3(new_n314), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n467), .A2(new_n472), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n316), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n500), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n497), .A2(new_n506), .A3(KEYINPUT84), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n320), .A2(new_n323), .A3(new_n233), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n300), .A2(new_n513), .A3(new_n233), .A4(G87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT22), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n233), .A2(G107), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT23), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT22), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n258), .A2(G116), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  XNOR2_X1  g0322(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(new_n523), .A3(new_n519), .A4(new_n517), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n347), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n518), .A2(new_n267), .A3(G13), .ZN(new_n529));
  XOR2_X1   g0329(.A(new_n529), .B(KEYINPUT25), .Z(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n210), .B2(new_n489), .ZN(new_n531));
  INV_X1    g0331(.A(G41), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT5), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n287), .A2(new_n534), .A3(new_n288), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT79), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n535), .A2(new_n536), .A3(new_n468), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n535), .B2(new_n468), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n292), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n215), .A2(new_n301), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n225), .A2(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n320), .A2(new_n541), .A3(new_n323), .A4(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G294), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n257), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n305), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n535), .A2(new_n468), .A3(new_n533), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(G264), .A3(new_n282), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n316), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n546), .A2(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n539), .ZN(new_n553));
  INV_X1    g0353(.A(G179), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n528), .A2(new_n531), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n509), .A2(new_n510), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G97), .A2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n211), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n560), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n209), .A2(KEYINPUT6), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n211), .A3(new_n563), .A4(new_n558), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n233), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n262), .A2(new_n206), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n338), .A2(G107), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n347), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n268), .A2(G97), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n489), .A2(new_n209), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n300), .A2(KEYINPUT4), .A3(G244), .A4(new_n301), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G283), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n336), .A2(new_n221), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(KEYINPUT4), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n300), .A2(G250), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n301), .B1(new_n577), .B2(KEYINPUT4), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n305), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n547), .A2(G257), .A3(new_n282), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n539), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n579), .A2(G190), .A3(new_n539), .A4(new_n580), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n572), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n316), .ZN(new_n585));
  INV_X1    g0385(.A(new_n570), .ZN(new_n586));
  INV_X1    g0386(.A(new_n571), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n210), .B1(new_n335), .B2(new_n337), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n588), .A2(new_n565), .A3(new_n566), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n587), .C1(new_n589), .C2(new_n347), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n579), .A2(new_n314), .A3(new_n539), .A4(new_n580), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n528), .A2(new_n531), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n540), .A2(G190), .A3(new_n549), .ZN(new_n595));
  AOI21_X1  g0395(.A(G200), .B1(new_n552), .B2(new_n539), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G264), .A2(G1698), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n300), .B(new_n600), .C1(new_n225), .C2(G1698), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n305), .C1(G303), .C2(new_n300), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n547), .A2(G270), .A3(new_n282), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n539), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n554), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n574), .B(new_n233), .C1(G33), .C2(new_n209), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G20), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n265), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G116), .B(new_n488), .C1(new_n388), .C2(new_n389), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n269), .A2(new_n607), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n604), .A2(new_n614), .A3(G169), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n604), .A2(G200), .ZN(new_n619));
  INV_X1    g0419(.A(new_n614), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n539), .A2(G190), .A3(new_n602), .A4(new_n603), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n604), .A2(new_n614), .A3(KEYINPUT21), .A4(G169), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n615), .A2(new_n618), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n593), .A2(new_n599), .A3(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n458), .A2(new_n557), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(new_n318), .ZN(new_n627));
  INV_X1    g0427(.A(new_n379), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n449), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n366), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n627), .B1(new_n631), .B2(new_n312), .ZN(new_n632));
  INV_X1    g0432(.A(new_n458), .ZN(new_n633));
  INV_X1    g0433(.A(new_n502), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT87), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n504), .A2(new_n635), .A3(new_n316), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT87), .B1(new_n492), .B2(G169), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n498), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT88), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n636), .A2(new_n637), .A3(new_n640), .A4(new_n498), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI211_X1 g0442(.A(new_n490), .B(new_n473), .C1(G190), .C2(new_n492), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n642), .A2(new_n592), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n592), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n509), .A2(new_n510), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n618), .A2(new_n615), .A3(new_n623), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n651), .B2(new_n556), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n597), .A2(new_n528), .A3(new_n531), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n584), .A2(new_n592), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n642), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n646), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n633), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n632), .A2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(new_n556), .ZN(new_n660));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G20), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n267), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT89), .ZN(new_n670));
  INV_X1    g0470(.A(new_n668), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n599), .B(new_n556), .C1(new_n594), .C2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n651), .A2(new_n668), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n660), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n614), .A2(new_n668), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n624), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n651), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n673), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(G399));
  NAND2_X1  g0485(.A1(new_n287), .A2(new_n288), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n236), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G1), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n480), .A2(G116), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n230), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n509), .A2(new_n645), .A3(new_n647), .A4(new_n510), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n644), .B2(new_n645), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n652), .A2(new_n655), .ZN(new_n697));
  INV_X1    g0497(.A(new_n642), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n671), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT92), .B(new_n671), .C1(new_n696), .C2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(KEYINPUT29), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n657), .A2(new_n671), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(new_n625), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n509), .A2(new_n510), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n556), .A4(new_n671), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n550), .A2(new_n313), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n504), .A3(new_n581), .A4(new_n604), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n492), .A2(new_n579), .A3(new_n539), .A4(new_n580), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT90), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT30), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(new_n552), .A3(new_n605), .A4(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n539), .A2(new_n603), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(G179), .A3(new_n552), .A4(new_n602), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n715), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n711), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n721), .B2(new_n668), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT91), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n668), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT91), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n722), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n709), .A2(new_n725), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n704), .A2(new_n706), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n694), .B1(new_n734), .B2(G1), .ZN(G364));
  NAND2_X1  g0535(.A1(new_n662), .A2(G45), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n690), .A2(G1), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n233), .A2(G190), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n313), .A2(new_n367), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n233), .A2(new_n369), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n313), .A2(new_n367), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n739), .A2(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G179), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n300), .B1(new_n748), .B2(G329), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n367), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n746), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n749), .B1(new_n750), .B2(new_n752), .C1(new_n544), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n742), .A2(new_n751), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n745), .B(new_n756), .C1(G303), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G326), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n314), .A2(new_n233), .A3(new_n367), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n765), .A2(G190), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n765), .A2(new_n369), .A3(new_n766), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  OAI221_X1 g0569(.A(new_n762), .B1(new_n763), .B2(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT96), .ZN(new_n771));
  INV_X1    g0571(.A(new_n767), .ZN(new_n772));
  INV_X1    g0572(.A(new_n768), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G50), .A2(new_n772), .B1(new_n773), .B2(G68), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n748), .A2(G159), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n760), .A2(new_n214), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n300), .B1(new_n752), .B2(new_n210), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n754), .A2(G97), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n741), .B2(new_n206), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n776), .A2(new_n777), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n774), .B(new_n781), .C1(new_n202), .C2(new_n743), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n232), .B1(G20), .B2(new_n316), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n738), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G13), .A2(G33), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n785), .B1(new_n681), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n788), .A2(new_n784), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n688), .A2(new_n300), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n231), .A2(new_n293), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(new_n251), .C2(new_n293), .ZN(new_n794));
  NAND3_X1  g0594(.A1(G355), .A2(new_n300), .A3(new_n236), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(G116), .C2(new_n236), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n790), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT97), .Z(new_n798));
  OR2_X1    g0598(.A1(new_n681), .A2(G330), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n682), .A3(new_n737), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(G396));
  NAND2_X1  g0601(.A1(new_n398), .A2(new_n668), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n401), .A2(new_n802), .B1(new_n404), .B2(new_n405), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n404), .A2(new_n405), .A3(new_n671), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n657), .A2(new_n671), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n401), .A2(new_n802), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n804), .B1(new_n809), .B2(new_n407), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n705), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n705), .A2(new_n810), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(KEYINPUT99), .B2(new_n807), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT100), .B1(new_n814), .B2(new_n732), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT100), .ZN(new_n816));
  INV_X1    g0616(.A(new_n732), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n817), .C1(new_n811), .C2(new_n813), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n814), .A2(new_n732), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n815), .A2(new_n737), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G303), .A2(new_n772), .B1(new_n773), .B2(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n607), .A2(new_n741), .B1(new_n743), .B2(new_n544), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n779), .B1(new_n214), .B2(new_n752), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n336), .B1(new_n747), .B2(new_n739), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n821), .B(new_n825), .C1(new_n210), .C2(new_n760), .ZN(new_n826));
  INV_X1    g0626(.A(G137), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n767), .B1(new_n768), .B2(new_n260), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  INV_X1    g0629(.A(G143), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n743), .C1(new_n340), .C2(new_n741), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n752), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G68), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n835), .C1(new_n202), .C2(new_n755), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n336), .B1(new_n748), .B2(G132), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n219), .B2(new_n760), .C1(new_n831), .C2(new_n832), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n826), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n738), .B1(new_n839), .B2(new_n784), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n784), .A2(new_n786), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(G77), .B2(new_n842), .C1(new_n787), .C2(new_n806), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n820), .A2(new_n843), .ZN(G384));
  NAND2_X1  g0644(.A1(new_n379), .A2(KEYINPUT101), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT101), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n375), .A2(new_n846), .A3(new_n378), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n845), .A2(new_n366), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n666), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n364), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n353), .A2(new_n850), .A3(new_n372), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n353), .A2(new_n850), .A3(new_n854), .A4(new_n372), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n848), .A2(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT102), .B1(new_n856), .B2(KEYINPUT38), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n375), .A2(new_n846), .A3(new_n378), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n846), .B1(new_n375), .B2(new_n378), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n850), .B1(new_n862), .B2(new_n366), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n853), .A2(new_n855), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n858), .B(new_n859), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n366), .A2(new_n379), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n851), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n857), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n438), .A2(new_n448), .A3(new_n671), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n868), .A2(new_n864), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n859), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n872), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n355), .A2(new_n365), .A3(new_n666), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n807), .A2(new_n804), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n869), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n438), .A2(new_n448), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n448), .A2(new_n668), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n457), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n448), .B(new_n668), .C1(new_n630), .C2(new_n438), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n878), .A2(new_n879), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n704), .A2(new_n706), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n633), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n632), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n888), .B(new_n891), .Z(new_n892));
  NOR3_X1   g0692(.A1(new_n557), .A2(new_n625), .A3(new_n668), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n728), .A2(new_n722), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n806), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n884), .B2(new_n885), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n870), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT40), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n723), .A2(new_n724), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n810), .B1(new_n709), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(KEYINPUT103), .A2(KEYINPUT40), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n886), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n881), .C1(new_n896), .C2(KEYINPUT103), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n709), .A2(new_n899), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n905), .A2(new_n449), .A3(new_n403), .A4(new_n457), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(G330), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n892), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n267), .B2(new_n662), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n561), .A2(new_n564), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n607), .B1(new_n911), .B2(KEYINPUT35), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n234), .C1(KEYINPUT35), .C2(new_n911), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n231), .A2(G77), .A3(new_n332), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n201), .A2(new_n203), .ZN(new_n916));
  OAI211_X1 g0716(.A(G1), .B(new_n661), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n914), .A3(new_n917), .ZN(G367));
  AOI211_X1 g0718(.A(new_n643), .B(new_n642), .C1(new_n490), .C2(new_n668), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT104), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n698), .A2(new_n495), .A3(new_n671), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n788), .ZN(new_n923));
  INV_X1    g0723(.A(new_n792), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n791), .B1(new_n236), .B2(new_n501), .C1(new_n247), .C2(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n544), .A2(new_n768), .B1(new_n767), .B2(new_n739), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n834), .A2(G97), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n210), .B2(new_n755), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n300), .B(new_n928), .C1(G317), .C2(new_n748), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT46), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n760), .B2(new_n607), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n761), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  INV_X1    g0732(.A(new_n741), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(G283), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n929), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n743), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n926), .B(new_n935), .C1(G303), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(G150), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n830), .A2(new_n767), .B1(new_n768), .B2(new_n340), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n754), .A2(G68), .ZN(new_n940));
  INV_X1    g0740(.A(new_n201), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n940), .B1(new_n827), .B2(new_n747), .C1(new_n941), .C2(new_n741), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n336), .B1(new_n834), .B2(G77), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT109), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n944), .B(new_n945), .C1(new_n202), .C2(new_n760), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n939), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n937), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n738), .B1(new_n950), .B2(new_n784), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n923), .A2(new_n925), .A3(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n736), .A2(G1), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n593), .B1(new_n572), .B2(new_n671), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n647), .A2(new_n668), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT44), .B1(new_n678), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  INV_X1    g0760(.A(new_n958), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n677), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n677), .B2(new_n961), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n677), .A2(new_n963), .A3(new_n961), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n959), .B(new_n962), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n684), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT108), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n959), .A2(new_n962), .ZN(new_n970));
  INV_X1    g0770(.A(new_n966), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n964), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n684), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n967), .A2(new_n968), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n673), .B(new_n674), .Z(new_n977));
  OR2_X1    g0777(.A1(new_n683), .A2(KEYINPUT107), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n733), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n975), .A2(new_n976), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n734), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n689), .B(KEYINPUT41), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n955), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT43), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n922), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n675), .A2(new_n956), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n592), .B1(new_n956), .B2(new_n556), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n671), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT106), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n922), .A2(new_n985), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT105), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n684), .A2(new_n961), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n994), .B(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n953), .B1(new_n984), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n980), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n690), .B1(new_n979), .B2(new_n733), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n752), .A2(new_n607), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n773), .A2(G311), .B1(G317), .B2(new_n936), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n744), .B2(new_n767), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G303), .B2(new_n933), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT48), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n760), .A2(new_n544), .B1(new_n750), .B2(new_n755), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT111), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n336), .B1(new_n763), .B2(new_n747), .C1(new_n1012), .C2(KEYINPUT49), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1005), .B(new_n1013), .C1(KEYINPUT49), .C2(new_n1012), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n340), .A2(new_n767), .B1(new_n768), .B2(new_n349), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n760), .A2(new_n206), .B1(new_n203), .B2(new_n741), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n743), .A2(new_n219), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n336), .B1(new_n748), .B2(G150), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n754), .A2(new_n394), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n927), .A3(new_n1019), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n784), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n738), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n256), .A2(new_n219), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n692), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n293), .C1(KEYINPUT50), .C2(new_n1024), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G68), .B2(G77), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n792), .B1(new_n244), .B2(new_n293), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n692), .A2(new_n236), .A3(new_n300), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n236), .A2(G107), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n791), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1022), .A2(new_n1023), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT112), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n673), .A2(new_n789), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1004), .B1(new_n955), .B2(new_n979), .C1(new_n1034), .C2(new_n1035), .ZN(G393));
  INV_X1    g0836(.A(new_n975), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n976), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n967), .A2(KEYINPUT113), .A3(new_n968), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT114), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT114), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n975), .A2(new_n1043), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n954), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1002), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1046), .A2(new_n689), .A3(new_n981), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n767), .A2(new_n260), .B1(new_n340), .B2(new_n743), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT51), .Z(new_n1049));
  OAI22_X1  g0849(.A1(new_n768), .A2(new_n941), .B1(new_n349), .B2(new_n741), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT115), .Z(new_n1051));
  NAND2_X1  g0851(.A1(new_n754), .A2(G77), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n300), .C1(new_n830), .C2(new_n747), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n760), .A2(new_n203), .B1(new_n214), .B2(new_n752), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n767), .A2(new_n1057), .B1(new_n739), .B2(new_n743), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT52), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n834), .A2(G107), .B1(new_n754), .B2(G116), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n300), .B1(new_n748), .B2(G322), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n544), .C2(new_n741), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n773), .B2(G303), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1060), .B(new_n1066), .C1(G283), .C2(new_n761), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n784), .B1(new_n1056), .B2(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n791), .B1(new_n209), .B2(new_n236), .C1(new_n254), .C2(new_n924), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n961), .A2(new_n788), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n1023), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1045), .A2(new_n1047), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT117), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1045), .A2(new_n1047), .A3(KEYINPUT117), .A4(new_n1071), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(G390));
  NAND2_X1  g0876(.A1(new_n872), .A2(new_n877), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n880), .A2(new_n886), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n873), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n886), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1081), .A2(new_n732), .A3(new_n810), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n702), .A2(new_n703), .A3(new_n804), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n803), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n886), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n870), .A2(new_n873), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1080), .A2(new_n1082), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G330), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1081), .A2(new_n1089), .A3(new_n895), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n633), .A2(KEYINPUT118), .A3(G330), .A4(new_n905), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT118), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n906), .B2(new_n1089), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n890), .A2(new_n1097), .A3(new_n632), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n731), .A2(G330), .A3(new_n806), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n886), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n880), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT119), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n905), .B2(G330), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(G330), .C1(new_n893), .C2(new_n894), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n806), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1081), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1083), .A2(new_n1084), .B1(new_n1099), .B2(new_n886), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT120), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1081), .B(new_n1109), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1098), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1093), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1101), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1098), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1113), .A2(new_n689), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1077), .A2(new_n786), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n761), .A2(G150), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  AOI22_X1  g0922(.A1(G132), .A2(new_n936), .B1(new_n933), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n336), .B1(new_n834), .B2(new_n201), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(new_n340), .C2(new_n755), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G128), .A2(new_n772), .B1(new_n773), .B2(G137), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1126), .B(new_n1127), .C1(new_n1128), .C2(new_n747), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G283), .A2(new_n772), .B1(new_n773), .B2(G107), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n300), .B1(new_n748), .B2(G294), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n835), .A3(new_n1052), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1132), .B(new_n777), .C1(G116), .C2(new_n936), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1130), .B(new_n1133), .C1(new_n209), .C2(new_n741), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n738), .B1(new_n1135), .B2(new_n784), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1119), .B(new_n1136), .C1(new_n256), .C2(new_n842), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1093), .B2(new_n954), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT121), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1118), .B1(new_n1141), .B2(new_n1142), .ZN(G378));
  XOR2_X1   g0943(.A(new_n319), .B(KEYINPUT55), .Z(new_n1144));
  NAND2_X1  g0944(.A1(new_n273), .A2(new_n849), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1144), .B(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1089), .B1(new_n898), .B2(new_n903), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n888), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n888), .A2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n888), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n904), .A2(G330), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1147), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n888), .A2(new_n1148), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1115), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n689), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT123), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(KEYINPUT123), .A3(new_n689), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1158), .A2(new_n954), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n257), .B(new_n532), .C1(new_n752), .C2(new_n340), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n761), .A2(new_n1122), .B1(G150), .B2(new_n754), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n827), .B2(new_n741), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G132), .B2(new_n773), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n936), .A2(G128), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n1128), .C2(new_n767), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1171), .B1(new_n1176), .B2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n748), .A2(G124), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(KEYINPUT59), .C2(new_n1176), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G116), .A2(new_n772), .B1(new_n773), .B2(G97), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n760), .A2(new_n206), .B1(new_n501), .B2(new_n741), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n687), .A2(new_n300), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n834), .A2(G58), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n748), .A2(G283), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n940), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1180), .B(new_n1186), .C1(new_n210), .C2(new_n743), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT58), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1179), .B(new_n1188), .C1(new_n1182), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n737), .B1(new_n1190), .B2(new_n784), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n201), .B2(new_n842), .C1(new_n1147), .C2(new_n787), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1170), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT122), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1170), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1169), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1114), .A2(new_n954), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G294), .A2(new_n772), .B1(new_n773), .B2(G116), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n300), .B1(new_n748), .B2(G303), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1203), .B(new_n1019), .C1(new_n206), .C2(new_n752), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n210), .A2(new_n741), .B1(new_n743), .B2(new_n750), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1202), .B(new_n1206), .C1(new_n209), .C2(new_n760), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G132), .A2(new_n772), .B1(new_n773), .B2(new_n1122), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n760), .A2(new_n340), .B1(new_n260), .B2(new_n741), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n336), .B1(new_n748), .B2(G128), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n1183), .C1(new_n219), .C2(new_n755), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1208), .B(new_n1212), .C1(new_n827), .C2(new_n743), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT124), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n738), .B1(new_n1215), .B2(new_n784), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(G68), .B2(new_n842), .C1(new_n886), .C2(new_n787), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1201), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1098), .A2(new_n1111), .A3(new_n1101), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(new_n983), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1219), .B1(new_n1222), .B2(new_n1112), .ZN(G381));
  AND2_X1   g1023(.A1(new_n1118), .A2(new_n1139), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1199), .A2(new_n1224), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G384), .A3(G381), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1074), .A2(new_n1000), .A3(new_n1075), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1227), .A2(G396), .A3(G393), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(G407));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1225), .ZN(G409));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1168), .A2(G378), .A3(new_n1197), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1164), .A2(new_n983), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1224), .B1(new_n1193), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(G213), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(G343), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT60), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1112), .B1(new_n1239), .B2(new_n1220), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1098), .A2(new_n1111), .A3(new_n1101), .A4(KEYINPUT60), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1241), .A2(new_n689), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1218), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT125), .B1(new_n1243), .B2(G384), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(G384), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1220), .A2(new_n1239), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(new_n689), .A3(new_n1116), .A4(new_n1241), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1219), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1244), .A2(new_n1245), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AND4_X1   g1053(.A1(new_n1231), .A2(new_n1235), .A3(new_n1238), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1237), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1231), .B1(new_n1255), .B2(new_n1253), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1249), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1261));
  AOI211_X1 g1061(.A(KEYINPUT125), .B(G384), .C1(new_n1247), .C2(new_n1219), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1263), .B2(new_n1245), .ZN(new_n1264));
  AND4_X1   g1064(.A1(new_n1260), .A2(new_n1244), .A3(new_n1245), .A4(new_n1251), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1259), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1260), .A3(new_n1245), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1252), .A2(KEYINPUT126), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(G2897), .A4(new_n1237), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1258), .B1(new_n1270), .B2(new_n1255), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT127), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n1258), .C1(new_n1270), .C2(new_n1255), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1257), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(G396), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1074), .A2(new_n1000), .A3(new_n1075), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1000), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G390), .A2(G387), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1227), .A3(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1275), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT63), .B1(new_n1270), .B2(new_n1255), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1255), .A2(new_n1253), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1287), .B(new_n1288), .C1(new_n1289), .C2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1284), .A2(new_n1290), .ZN(G405));
  NAND2_X1  g1091(.A1(G375), .A2(new_n1224), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1283), .A2(new_n1232), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1283), .B1(new_n1232), .B2(new_n1292), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1252), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1232), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1288), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(new_n1253), .A3(new_n1293), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1299), .ZN(G402));
endmodule


