//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n202), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n215), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n207), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n248), .A2(new_n249), .B1(new_n207), .B2(G68), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n207), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n202), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n247), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT71), .Z(new_n255));
  OR2_X1    g0055(.A1(new_n255), .A2(KEYINPUT11), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n240), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n255), .A2(KEYINPUT11), .ZN(new_n261));
  OAI21_X1  g0061(.A(KEYINPUT68), .B1(new_n258), .B2(new_n247), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n257), .A2(new_n263), .A3(new_n215), .A4(new_n246), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(new_n206), .B2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G68), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n256), .A2(new_n260), .A3(new_n261), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT14), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  OAI21_X1  g0074(.A(G238), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n274), .B2(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G97), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n228), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G226), .B2(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n206), .A2(G274), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT64), .B(G45), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(G41), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n276), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n276), .A2(new_n291), .A3(KEYINPUT13), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n269), .B(G169), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n269), .B1(new_n297), .B2(G169), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n268), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n294), .A2(new_n295), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n268), .B1(new_n302), .B2(G190), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n297), .A2(G200), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(G77), .ZN(new_n308));
  INV_X1    g0108(.A(new_n247), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT8), .B(G58), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n252), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G20), .B2(G77), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  OR3_X1    g0113(.A1(new_n313), .A2(KEYINPUT67), .A3(new_n248), .ZN(new_n314));
  OAI21_X1  g0114(.A(KEYINPUT67), .B1(new_n313), .B2(new_n248), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n308), .B1(G77), .B2(new_n257), .C1(new_n309), .C2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT3), .B(G33), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(G238), .A3(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(G1698), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(G232), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G107), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n319), .B(new_n321), .C1(new_n322), .C2(new_n318), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n285), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT64), .A2(G45), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT64), .A2(G45), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G41), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n287), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n273), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(G244), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n317), .B1(G200), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(new_n298), .A3(new_n331), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n317), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G58), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n341), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT65), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n310), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n251), .A2(G20), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G20), .A2(G33), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n309), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n257), .A2(G50), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n247), .B1(new_n206), .B2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(G50), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n329), .B1(G226), .B2(new_n330), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G222), .A2(G1698), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n320), .A2(G223), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n318), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n285), .C1(G77), .C2(new_n318), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n336), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n298), .A3(new_n360), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n355), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XOR2_X1   g0164(.A(new_n364), .B(KEYINPUT66), .Z(new_n365));
  NOR2_X1   g0165(.A1(new_n340), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT18), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n281), .B2(G33), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n251), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n282), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(new_n318), .B2(G20), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n240), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n341), .A2(new_n240), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n347), .A2(KEYINPUT73), .A3(G159), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT73), .B1(new_n347), .B2(G159), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n368), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n318), .A2(new_n373), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n283), .B2(new_n207), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(KEYINPUT72), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n377), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n240), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n380), .B(KEYINPUT16), .C1(new_n381), .C2(new_n382), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n384), .B(new_n247), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n344), .A2(new_n257), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n344), .B2(new_n351), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OR2_X1    g0195(.A1(G223), .A2(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G226), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G1698), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n280), .A2(new_n396), .A3(new_n282), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n271), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n405), .B2(new_n329), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n290), .A2(KEYINPUT75), .A3(new_n404), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n290), .A2(new_n404), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n336), .B1(new_n409), .B2(new_n401), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n367), .B1(new_n395), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(KEYINPUT18), .B(new_n411), .C1(new_n392), .C2(new_n394), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n401), .A2(G190), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(new_n406), .A3(new_n407), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n409), .B2(new_n401), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n392), .A2(new_n394), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n394), .ZN(new_n425));
  OAI211_X1 g0225(.A(KEYINPUT72), .B(new_n376), .C1(new_n318), .C2(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n283), .A2(new_n374), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n283), .A2(new_n207), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT72), .B1(new_n429), .B2(new_n376), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n391), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n309), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n433), .B2(new_n384), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n416), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT10), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n361), .A2(new_n334), .B1(KEYINPUT69), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n439), .B1(G200), .B2(new_n361), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n354), .A2(KEYINPUT9), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(KEYINPUT69), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n445), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n307), .A2(new_n366), .A3(new_n437), .A4(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(G1698), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(new_n320), .ZN(new_n453));
  INV_X1    g0253(.A(G294), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n251), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n285), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n206), .A2(G45), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT5), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(G41), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n328), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT76), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n458), .B2(G41), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n459), .A2(G274), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G45), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(G41), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(new_n460), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(G264), .A3(new_n271), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n336), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n456), .A2(new_n298), .A3(new_n463), .A4(new_n468), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n280), .A2(new_n282), .A3(new_n207), .A4(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n318), .A2(new_n475), .A3(new_n207), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n207), .B2(G107), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n322), .A2(KEYINPUT23), .A3(G20), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n477), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n478), .B1(new_n477), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n247), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n309), .B(new_n257), .C1(G1), .C2(new_n251), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n258), .A2(new_n322), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  AOI22_X1  g0294(.A1(G107), .A2(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n472), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n456), .A2(G190), .A3(new_n463), .A4(new_n468), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n469), .A2(G200), .ZN(new_n498));
  AND4_X1   g0298(.A1(new_n487), .A2(new_n495), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT84), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(new_n470), .A3(new_n471), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT84), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n487), .A2(new_n495), .A3(new_n498), .A4(new_n497), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G283), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(new_n320), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n509), .A2(new_n510), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n285), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n467), .A2(G257), .A3(new_n271), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n514), .A2(new_n463), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT77), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT77), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(G200), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT78), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT78), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(G190), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n375), .A2(new_n377), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G97), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n528), .A2(new_n530), .A3(G107), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(G20), .B1(G77), .B2(new_n347), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n309), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n257), .A2(G97), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n488), .B2(new_n530), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n520), .A2(new_n524), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT78), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT78), .B1(new_n513), .B2(new_n515), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n336), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n513), .A2(new_n515), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n531), .B1(new_n528), .B2(new_n527), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n545), .A2(new_n207), .B1(new_n249), .B2(new_n252), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n322), .B1(new_n375), .B2(new_n377), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n247), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n538), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n544), .A2(new_n298), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n540), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n206), .B2(G33), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n262), .A2(new_n264), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G13), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(G1), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(G20), .A3(new_n553), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n246), .A2(new_n215), .B1(G20), .B2(new_n553), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n508), .B(new_n207), .C1(G33), .C2(new_n530), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n280), .A2(new_n282), .A3(G264), .A4(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(new_n320), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n318), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n285), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n467), .A2(G270), .A3(new_n271), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n463), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n563), .B1(new_n570), .B2(G200), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n334), .B2(new_n570), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n563), .A3(G169), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n569), .A2(new_n463), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n563), .A2(G179), .A3(new_n568), .A4(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n570), .A2(new_n563), .A3(KEYINPUT21), .A4(G169), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n572), .A2(new_n575), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n280), .A2(new_n282), .A3(new_n207), .A4(G68), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT81), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n345), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n318), .A2(KEYINPUT81), .A3(new_n207), .A4(G68), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n207), .B1(new_n277), .B2(new_n583), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G97), .A2(G107), .ZN(new_n589));
  INV_X1    g0389(.A(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n587), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n247), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n313), .A2(new_n258), .ZN(new_n596));
  OR2_X1    g0396(.A1(new_n488), .A2(new_n313), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT79), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n457), .A2(G250), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n285), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n271), .A2(KEYINPUT79), .A3(G250), .A4(new_n457), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n601), .A2(new_n602), .B1(G45), .B2(new_n288), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n280), .A2(new_n282), .A3(G238), .A4(new_n320), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n479), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n285), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n336), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n603), .A2(new_n607), .A3(new_n298), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n598), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(new_n607), .A3(G190), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT82), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n584), .B(new_n585), .C1(new_n592), .C2(new_n593), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(new_n247), .B1(new_n258), .B2(new_n313), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(G200), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n489), .A2(G87), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n611), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n552), .A2(new_n579), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n451), .A2(new_n506), .A3(new_n620), .ZN(G372));
  INV_X1    g0421(.A(new_n305), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n301), .B1(new_n622), .B2(new_n339), .ZN(new_n623));
  INV_X1    g0423(.A(new_n436), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n415), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n365), .B1(new_n626), .B2(new_n449), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n595), .A2(new_n596), .A3(new_n617), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n419), .B1(new_n603), .B2(new_n607), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT85), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT82), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n612), .B(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n615), .A2(new_n616), .A3(new_n633), .A4(new_n617), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n535), .A2(new_n538), .B1(new_n516), .B2(G179), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n522), .A2(new_n523), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n336), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n635), .A2(new_n638), .A3(new_n639), .A4(new_n611), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT26), .B1(new_n619), .B2(new_n551), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n611), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n504), .B1(new_n496), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n552), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n635), .A2(new_n611), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n642), .A2(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT86), .A4(new_n611), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n627), .B1(new_n450), .B2(new_n650), .ZN(G369));
  INV_X1    g0451(.A(new_n557), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT87), .B1(new_n652), .B2(G20), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT27), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n557), .A2(new_n655), .A3(new_n207), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n653), .B2(new_n656), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n501), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g0464(.A(new_n664), .B(KEYINPUT88), .Z(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n506), .ZN(new_n666));
  INV_X1    g0466(.A(new_n663), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n502), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n663), .A2(new_n563), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n644), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n579), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n666), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n663), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n676), .A2(new_n678), .B1(new_n496), .B2(new_n667), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n210), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n589), .A2(new_n590), .A3(new_n553), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT89), .Z(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(new_n684), .A3(new_n206), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n214), .B2(new_n682), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT90), .Z(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  INV_X1    g0488(.A(G330), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n540), .A2(new_n551), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n579), .A2(new_n619), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n506), .A2(new_n690), .A3(new_n691), .A4(new_n667), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT93), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n620), .A2(new_n694), .A3(new_n506), .A4(new_n667), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n603), .B2(new_n607), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n516), .A2(new_n697), .A3(new_n469), .A4(new_n570), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n570), .A2(new_n298), .ZN(new_n700));
  AND4_X1   g0500(.A1(new_n468), .A2(new_n456), .A3(new_n603), .A4(new_n607), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n522), .A2(new_n700), .A3(new_n523), .A4(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n541), .A2(new_n542), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n700), .A4(new_n701), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n667), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT92), .B1(new_n707), .B2(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n706), .A2(new_n709), .A3(new_n698), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n663), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT92), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT91), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n707), .A2(new_n717), .A3(KEYINPUT31), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n708), .A2(new_n714), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n689), .B1(new_n696), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n499), .B1(new_n677), .B2(new_n502), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n647), .A2(new_n690), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n635), .A2(new_n611), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT26), .B1(new_n725), .B2(new_n551), .ZN(new_n726));
  INV_X1    g0526(.A(new_n611), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n619), .A2(new_n551), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n639), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n722), .B1(new_n730), .B2(new_n667), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n663), .B1(new_n648), .B2(new_n649), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n721), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n688), .B1(new_n735), .B2(G1), .ZN(G364));
  NOR2_X1   g0536(.A1(new_n556), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n206), .B1(new_n737), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n682), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n210), .A2(G355), .A3(new_n318), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(new_n318), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n213), .B2(new_n289), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n244), .A2(new_n464), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(G116), .B2(new_n210), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n215), .B1(G20), .B2(new_n336), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n741), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n207), .A2(new_n334), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n298), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT96), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G58), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n419), .A2(G179), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n207), .A2(G190), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n283), .B1(new_n768), .B2(G107), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n756), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n755), .A2(new_n765), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n769), .B1(new_n249), .B2(new_n770), .C1(new_n590), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G159), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n207), .B1(new_n773), .B2(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n334), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n779), .A2(G97), .B1(G50), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n240), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n772), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n775), .A2(G329), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n787), .B1(new_n566), .B2(new_n771), .C1(new_n788), .C2(new_n770), .ZN(new_n789));
  INV_X1    g0589(.A(new_n761), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G322), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n283), .B1(new_n767), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI22_X1  g0594(.A1(new_n784), .A2(new_n794), .B1(new_n454), .B2(new_n778), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G326), .C2(new_n781), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n764), .A2(new_n786), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n750), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n754), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT97), .ZN(new_n800));
  INV_X1    g0600(.A(new_n749), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n672), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n672), .A2(G330), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n673), .A2(new_n741), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(G396));
  NOR2_X1   g0605(.A1(new_n750), .A2(new_n747), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n741), .B1(new_n249), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n768), .A2(G87), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n553), .B2(new_n770), .C1(new_n788), .C2(new_n774), .ZN(new_n809));
  INV_X1    g0609(.A(new_n771), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n318), .B1(new_n810), .B2(G107), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n783), .A2(G283), .B1(new_n781), .B2(G303), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(new_n530), .C2(new_n778), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n809), .B(new_n813), .C1(G294), .C2(new_n790), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  INV_X1    g0615(.A(new_n770), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G159), .B1(G137), .B2(new_n781), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n784), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n763), .B2(G143), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n283), .B1(new_n810), .B2(G50), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n779), .A2(G58), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n768), .A2(G68), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n775), .A2(G132), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n820), .B2(KEYINPUT34), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n815), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n317), .A2(new_n663), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n335), .A2(new_n339), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n317), .A2(new_n337), .A3(new_n338), .A4(new_n663), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT99), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n807), .B1(new_n798), .B2(new_n828), .C1(new_n833), .C2(new_n748), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n732), .B(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n721), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n721), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n741), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(G384));
  OR2_X1    g0640(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(G116), .A3(new_n216), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  XNOR2_X1  g0644(.A(new_n239), .B(KEYINPUT101), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n214), .B(G77), .C1(new_n341), .C2(new_n240), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n206), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n368), .B1(new_n390), .B2(new_n383), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n433), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n394), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n660), .B(new_n851), .C1(new_n416), .C2(new_n436), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n411), .A2(new_n661), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n851), .A2(new_n853), .B1(new_n434), .B2(new_n421), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n395), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n422), .A2(new_n855), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n852), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT105), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT17), .B1(new_n434), .B2(new_n421), .ZN(new_n866));
  AND4_X1   g0666(.A1(KEYINPUT17), .A2(new_n392), .A3(new_n394), .A4(new_n421), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n424), .A2(new_n435), .A3(KEYINPUT105), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n415), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n434), .A2(new_n661), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n870), .A2(KEYINPUT106), .A3(new_n871), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  OR3_X1    g0676(.A1(new_n856), .A2(new_n857), .A3(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n422), .A2(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n422), .A2(KEYINPUT103), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(KEYINPUT37), .C1(new_n856), .C2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n856), .B2(new_n857), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(new_n875), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n884));
  AOI21_X1  g0684(.A(new_n864), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n863), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n301), .A2(new_n663), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n339), .A2(new_n663), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n732), .B2(new_n833), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n861), .A2(new_n862), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n268), .A2(new_n663), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n306), .B(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n416), .A2(new_n661), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n890), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n733), .A2(new_n450), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n901), .A2(new_n627), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n883), .A2(new_n884), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n862), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n306), .A2(new_n896), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n895), .B1(new_n301), .B2(new_n305), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n833), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n711), .A2(new_n713), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n715), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n693), .B2(new_n695), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n861), .B2(new_n862), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n911), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n451), .A3(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n913), .A2(KEYINPUT40), .B1(new_n912), .B2(new_n915), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n450), .B2(new_n911), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(G330), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n903), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n206), .B2(new_n737), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n903), .A2(new_n922), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n848), .B1(new_n924), .B2(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n663), .A2(new_n628), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n647), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n611), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n540), .B(new_n551), .C1(new_n539), .C2(new_n667), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT107), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(new_n551), .C2(new_n667), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n496), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n663), .B1(new_n937), .B2(new_n551), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n676), .A3(new_n678), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n930), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT109), .Z(new_n942));
  NOR2_X1   g0742(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n936), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n675), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n679), .A2(new_n935), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT45), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n679), .A2(new_n935), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n675), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n676), .A2(new_n678), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n668), .A2(new_n678), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(KEYINPUT110), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(new_n673), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n734), .B1(new_n954), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n682), .B(KEYINPUT41), .Z(new_n963));
  OAI21_X1  g0763(.A(new_n738), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n944), .A2(new_n674), .A3(new_n936), .A4(new_n945), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n948), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n753), .B1(new_n210), .B2(new_n313), .ZN(new_n967));
  INV_X1    g0767(.A(new_n743), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n234), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n740), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n763), .A2(G303), .B1(G311), .B2(new_n781), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n767), .A2(new_n530), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n318), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT112), .B(G317), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n975), .B1(new_n792), .B2(new_n770), .C1(new_n774), .C2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n771), .A2(new_n553), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n784), .A2(new_n454), .B1(new_n778), .B2(new_n322), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n972), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n790), .A2(G150), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n318), .B1(new_n767), .B2(new_n249), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G159), .B2(new_n783), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n778), .A2(new_n240), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n781), .B2(G143), .ZN(new_n987));
  INV_X1    g0787(.A(G137), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n771), .A2(new_n341), .B1(new_n774), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G50), .B2(new_n816), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n983), .A2(new_n985), .A3(new_n987), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n970), .B1(new_n993), .B2(new_n750), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n801), .B2(new_n929), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT113), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n966), .A2(new_n996), .ZN(G387));
  NAND3_X1  g0797(.A1(new_n684), .A2(new_n210), .A3(new_n318), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(G107), .B2(new_n210), .ZN(new_n999));
  AOI211_X1 g0799(.A(G45), .B(new_n684), .C1(G68), .C2(G77), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n310), .A2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT50), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n968), .B1(new_n231), .B2(new_n289), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n999), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G77), .A2(new_n810), .B1(new_n775), .B2(G150), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n240), .B2(new_n770), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n778), .A2(new_n313), .ZN(new_n1011));
  NOR4_X1   g0811(.A1(new_n1010), .A2(new_n283), .A3(new_n974), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n781), .A2(G159), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT115), .Z(new_n1014));
  AOI22_X1  g0814(.A1(new_n790), .A2(G50), .B1(new_n344), .B2(new_n783), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n816), .A2(G303), .B1(G322), .B2(new_n781), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n788), .B2(new_n784), .C1(new_n762), .C2(new_n976), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n810), .A2(G294), .B1(new_n779), .B2(G283), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT49), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n767), .A2(new_n553), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n318), .B(new_n1025), .C1(G326), .C2(new_n775), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1016), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n740), .B1(new_n752), .B2(new_n1008), .C1(new_n1027), .C2(new_n798), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT116), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1028), .A2(new_n1029), .B1(new_n668), .B2(new_n801), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n739), .B2(new_n961), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n960), .A2(new_n734), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n682), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n735), .B2(new_n961), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n1034), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n954), .B2(new_n1033), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1033), .B2(new_n954), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n947), .A2(new_n749), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n753), .B1(new_n530), .B2(new_n210), .C1(new_n238), .C2(new_n968), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT118), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n740), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(G159), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n781), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n761), .A2(new_n1045), .B1(new_n818), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n775), .A2(G143), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n240), .B2(new_n771), .C1(new_n310), .C2(new_n770), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n778), .A2(new_n249), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n808), .B(new_n318), .C1(new_n202), .C2(new_n784), .ZN(new_n1052));
  OR4_X1    g0852(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n790), .A2(G311), .B1(G317), .B2(new_n781), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n283), .B1(new_n767), .B2(new_n322), .C1(new_n784), .C2(new_n566), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G294), .A2(new_n816), .B1(new_n775), .B2(G322), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n792), .B2(new_n771), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1056), .B(new_n1058), .C1(G116), .C2(new_n779), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n798), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1044), .B(new_n1061), .C1(new_n1043), .C2(new_n1042), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n954), .A2(new_n739), .B1(new_n1041), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1040), .A2(new_n1063), .ZN(G390));
  NOR2_X1   g0864(.A1(new_n906), .A2(new_n907), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n888), .B1(new_n892), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n886), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n720), .A2(new_n833), .A3(new_n897), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n730), .A2(new_n833), .A3(new_n667), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n891), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n889), .B1(new_n1071), .B2(new_n897), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT119), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n905), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n905), .B2(new_n1072), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1067), .B(new_n1068), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n918), .A2(new_n451), .A3(G330), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n627), .B(new_n1077), .C1(new_n450), .C2(new_n733), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n897), .B1(new_n720), .B2(new_n833), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n908), .A2(new_n911), .A3(new_n689), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n893), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n833), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n911), .A2(new_n689), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1068), .B(new_n1082), .C1(new_n1084), .C2(new_n897), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1078), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n888), .B1(new_n1082), .B2(new_n1065), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT119), .B1(new_n1087), .B2(new_n885), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n905), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1088), .A2(new_n1089), .B1(new_n886), .B2(new_n1066), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1080), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1076), .B(new_n1086), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(KEYINPUT120), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1067), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1080), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT120), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n1076), .A4(new_n1086), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1076), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1086), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1034), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(new_n739), .A3(new_n1076), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n806), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n740), .B1(new_n344), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n824), .B1(new_n530), .B2(new_n770), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G294), .B2(new_n775), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n790), .A2(G116), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n318), .B(new_n1051), .C1(G87), .C2(new_n810), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n783), .A2(G107), .B1(new_n781), .B2(G283), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n784), .A2(new_n988), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n318), .B1(new_n774), .B2(new_n1113), .C1(new_n202), .C2(new_n767), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n771), .A2(new_n818), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1112), .B(new_n1114), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(G132), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT54), .B(G143), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT121), .Z(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1118), .B1(new_n1119), .B2(new_n761), .C1(new_n770), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n781), .A2(G128), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n1045), .B2(new_n778), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1111), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT123), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n798), .B1(new_n1126), .B2(KEYINPUT123), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1105), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n887), .B2(new_n748), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1103), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1102), .A2(new_n1131), .ZN(G378));
  NAND3_X1  g0932(.A1(new_n890), .A2(new_n898), .A3(new_n899), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n449), .A2(new_n364), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n661), .A2(new_n354), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1134), .B(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n917), .B2(G330), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n920), .A2(new_n689), .A3(new_n1141), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1133), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n917), .A2(G330), .A3(new_n1142), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1141), .B1(new_n920), .B2(new_n689), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n900), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1141), .A2(new_n747), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n283), .A2(new_n328), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G283), .B2(new_n775), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n313), .B2(new_n770), .C1(new_n761), .C2(new_n322), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n771), .A2(new_n249), .B1(new_n767), .B2(new_n341), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n784), .A2(new_n530), .B1(new_n1046), .B2(new_n553), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1153), .A2(new_n986), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1151), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1122), .A2(new_n771), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT124), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n770), .A2(new_n988), .B1(new_n778), .B2(new_n818), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n784), .A2(new_n1119), .B1(new_n1046), .B2(new_n1113), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n790), .C2(G128), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1162), .A2(KEYINPUT124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n251), .B(new_n328), .C1(new_n767), .C2(new_n1045), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G124), .C2(new_n775), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1160), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(new_n798), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n741), .B(new_n1174), .C1(new_n202), .C2(new_n806), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1149), .A2(new_n739), .B1(new_n1150), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1078), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1098), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1034), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1078), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1149), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1177), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  INV_X1    g0987(.A(new_n963), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1081), .A2(new_n1085), .A3(new_n1078), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1100), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n738), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1065), .A2(new_n747), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n740), .B1(G68), .B2(new_n1104), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT125), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n790), .A2(G283), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n318), .B(new_n1011), .C1(G77), .C2(new_n768), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n783), .A2(G116), .B1(new_n781), .B2(G294), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n771), .A2(new_n530), .B1(new_n770), .B2(new_n322), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G303), .B2(new_n775), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n762), .A2(new_n988), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1121), .A2(new_n783), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n771), .A2(new_n1045), .B1(new_n770), .B2(new_n818), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G128), .B2(new_n775), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n781), .A2(G132), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n318), .B1(new_n767), .B2(new_n341), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G50), .B2(new_n779), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1200), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1194), .B1(new_n1209), .B2(new_n750), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1191), .B1(new_n1192), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1190), .A2(new_n1211), .ZN(G381));
  OR2_X1    g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1213), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n966), .A2(new_n996), .ZN(new_n1215));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1186), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n662), .A2(G213), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1186), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  NAND3_X1  g1021(.A1(new_n1179), .A2(new_n1188), .A3(new_n1149), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G378), .B1(new_n1222), .B2(new_n1176), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1186), .B2(G378), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT127), .B1(new_n1224), .B2(new_n1219), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1189), .B1(new_n1086), .B2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1081), .A2(new_n1085), .A3(new_n1078), .A4(KEYINPUT60), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n682), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1211), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(G384), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1222), .A2(new_n1176), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1216), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1149), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1149), .A2(KEYINPUT57), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n682), .B1(new_n1235), .B2(new_n1183), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1176), .C1(new_n1234), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT127), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1218), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1225), .A2(new_n1231), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT62), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1218), .A3(new_n1231), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(KEYINPUT126), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1238), .A2(new_n1231), .A3(new_n1247), .A4(new_n1218), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1219), .A2(G2897), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1231), .B(new_n1250), .Z(new_n1251));
  AOI21_X1  g1051(.A(new_n1239), .B1(new_n1238), .B2(new_n1218), .ZN(new_n1252));
  AOI211_X1 g1052(.A(KEYINPUT127), .B(new_n1219), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1242), .A2(new_n1243), .A3(new_n1249), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G390), .B1(new_n1213), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1213), .A2(G390), .A3(new_n1256), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n966), .A3(new_n996), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  OAI21_X1  g1061(.A(G387), .B1(new_n1261), .B2(new_n1257), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1255), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1238), .A2(new_n1218), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1265), .A2(new_n1251), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1263), .A2(new_n1266), .A3(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1267), .B(new_n1270), .C1(new_n1269), .C2(new_n1241), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1264), .A2(new_n1271), .ZN(G405));
  XNOR2_X1  g1072(.A(new_n1186), .B(G378), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1273), .A2(new_n1231), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1231), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(new_n1263), .Z(G402));
endmodule


