

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746;

  OR2_X1 U365 ( .A1(n393), .A2(n390), .ZN(n677) );
  NOR2_X1 U366 ( .A1(n636), .A2(n707), .ZN(n511) );
  OR2_X1 U367 ( .A1(n719), .A2(G902), .ZN(n467) );
  NAND2_X1 U368 ( .A1(n494), .A2(n493), .ZN(n377) );
  NOR2_X2 U369 ( .A1(n423), .A2(n420), .ZN(n448) );
  NAND2_X1 U370 ( .A1(n582), .A2(n584), .ZN(n657) );
  INV_X1 U371 ( .A(G143), .ZN(n489) );
  XNOR2_X1 U372 ( .A(G104), .B(G110), .ZN(n461) );
  INV_X2 U373 ( .A(n377), .ZN(n365) );
  NAND2_X1 U374 ( .A1(n401), .A2(n350), .ZN(n733) );
  NOR2_X1 U375 ( .A1(n407), .A2(n404), .ZN(n589) );
  XNOR2_X1 U376 ( .A(n465), .B(n463), .ZN(n742) );
  NOR2_X1 U377 ( .A1(n612), .A2(n611), .ZN(n624) );
  XNOR2_X1 U378 ( .A(n605), .B(n604), .ZN(n612) );
  XNOR2_X1 U379 ( .A(n677), .B(n484), .ZN(n622) );
  XNOR2_X1 U380 ( .A(n538), .B(n537), .ZN(n566) );
  XNOR2_X1 U381 ( .A(n476), .B(n473), .ZN(n547) );
  XNOR2_X1 U382 ( .A(n501), .B(n488), .ZN(n529) );
  XNOR2_X1 U383 ( .A(n461), .B(G107), .ZN(n419) );
  XNOR2_X1 U384 ( .A(G119), .B(G101), .ZN(n389) );
  XNOR2_X1 U385 ( .A(G116), .B(KEYINPUT88), .ZN(n388) );
  NAND2_X1 U386 ( .A1(n342), .A2(n343), .ZN(n705) );
  AND2_X1 U387 ( .A1(n669), .A2(n668), .ZN(n342) );
  NOR2_X1 U388 ( .A1(n703), .A2(G953), .ZN(n343) );
  XNOR2_X1 U389 ( .A(n387), .B(n462), .ZN(n366) );
  XNOR2_X1 U390 ( .A(n428), .B(n447), .ZN(n367) );
  XNOR2_X1 U391 ( .A(n508), .B(n507), .ZN(n707) );
  XNOR2_X2 U392 ( .A(n399), .B(n452), .ZN(n711) );
  XNOR2_X1 U393 ( .A(n441), .B(n399), .ZN(n559) );
  XNOR2_X1 U394 ( .A(n566), .B(n565), .ZN(n585) );
  NAND2_X1 U395 ( .A1(n398), .A2(n622), .ZN(n483) );
  NAND2_X1 U396 ( .A1(n742), .A2(n647), .ZN(n621) );
  NAND2_X1 U397 ( .A1(n635), .A2(n634), .ZN(n426) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n499) );
  NOR2_X2 U399 ( .A1(n397), .A2(n673), .ZN(n615) );
  NAND2_X1 U400 ( .A1(n469), .A2(n468), .ZN(n493) );
  INV_X1 U401 ( .A(KEYINPUT2), .ZN(n468) );
  XNOR2_X1 U402 ( .A(n567), .B(KEYINPUT41), .ZN(n684) );
  NAND2_X1 U403 ( .A1(n395), .A2(n394), .ZN(n393) );
  NOR2_X1 U404 ( .A1(n559), .A2(n391), .ZN(n390) );
  NAND2_X1 U405 ( .A1(G472), .A2(G902), .ZN(n394) );
  INV_X1 U406 ( .A(KEYINPUT47), .ZN(n406) );
  INV_X1 U407 ( .A(KEYINPUT81), .ZN(n431) );
  XNOR2_X1 U408 ( .A(n359), .B(G125), .ZN(n514) );
  INV_X1 U409 ( .A(G146), .ZN(n359) );
  XNOR2_X1 U410 ( .A(G902), .B(KEYINPUT15), .ZN(n552) );
  OR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n561) );
  XNOR2_X1 U412 ( .A(G143), .B(G122), .ZN(n516) );
  XOR2_X1 U413 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n517) );
  XNOR2_X1 U414 ( .A(G113), .B(G104), .ZN(n522) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n523) );
  XNOR2_X1 U416 ( .A(n580), .B(KEYINPUT46), .ZN(n383) );
  XNOR2_X1 U417 ( .A(n595), .B(KEYINPUT48), .ZN(n596) );
  INV_X1 U418 ( .A(KEYINPUT68), .ZN(n595) );
  NAND2_X1 U419 ( .A1(n621), .A2(KEYINPUT44), .ZN(n425) );
  NOR2_X1 U420 ( .A1(n744), .A2(KEYINPUT84), .ZN(n424) );
  XNOR2_X1 U421 ( .A(n514), .B(KEYINPUT10), .ZN(n544) );
  NOR2_X1 U422 ( .A1(n716), .A2(G902), .ZN(n538) );
  XNOR2_X1 U423 ( .A(n498), .B(n349), .ZN(n441) );
  XOR2_X1 U424 ( .A(KEYINPUT8), .B(n532), .Z(n549) );
  NAND2_X1 U425 ( .A1(G234), .A2(n704), .ZN(n532) );
  INV_X1 U426 ( .A(G134), .ZN(n488) );
  XNOR2_X1 U427 ( .A(n492), .B(n451), .ZN(n450) );
  XNOR2_X1 U428 ( .A(n536), .B(KEYINPUT9), .ZN(n451) );
  XNOR2_X1 U429 ( .A(G122), .B(KEYINPUT101), .ZN(n533) );
  INV_X1 U430 ( .A(n351), .ZN(n376) );
  NAND2_X1 U431 ( .A1(n381), .A2(n379), .ZN(n378) );
  NOR2_X1 U432 ( .A1(n380), .A2(n721), .ZN(n379) );
  NOR2_X1 U433 ( .A1(n351), .A2(G475), .ZN(n380) );
  XNOR2_X1 U434 ( .A(n728), .B(n346), .ZN(n508) );
  XNOR2_X1 U435 ( .A(n579), .B(n578), .ZN(n597) );
  NOR2_X1 U436 ( .A1(n576), .A2(n586), .ZN(n579) );
  NOR2_X1 U437 ( .A1(n630), .A2(n444), .ZN(n605) );
  XNOR2_X1 U438 ( .A(n446), .B(n445), .ZN(n444) );
  INV_X1 U439 ( .A(KEYINPUT64), .ZN(n464) );
  NAND2_X1 U440 ( .A1(n411), .A2(KEYINPUT28), .ZN(n410) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n555) );
  XNOR2_X1 U442 ( .A(n527), .B(n526), .ZN(n584) );
  INV_X1 U443 ( .A(KEYINPUT6), .ZN(n484) );
  NAND2_X1 U444 ( .A1(n378), .A2(n356), .ZN(n375) );
  INV_X1 U445 ( .A(n378), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n455), .B(n453), .ZN(n452) );
  XNOR2_X1 U447 ( .A(n515), .B(n454), .ZN(n453) );
  AND2_X1 U448 ( .A1(n493), .A2(G210), .ZN(n362) );
  AND2_X1 U449 ( .A1(n632), .A2(n405), .ZN(n404) );
  XNOR2_X1 U450 ( .A(n408), .B(n431), .ZN(n407) );
  XNOR2_X1 U451 ( .A(n495), .B(KEYINPUT67), .ZN(n502) );
  INV_X1 U452 ( .A(KEYINPUT4), .ZN(n495) );
  XNOR2_X1 U453 ( .A(n438), .B(n437), .ZN(n691) );
  INV_X1 U454 ( .A(KEYINPUT104), .ZN(n437) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(G131), .Z(n497) );
  XNOR2_X1 U456 ( .A(G116), .B(G107), .ZN(n528) );
  XOR2_X1 U457 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n534) );
  AND2_X1 U458 ( .A1(n493), .A2(n353), .ZN(n363) );
  XNOR2_X1 U459 ( .A(n529), .B(n486), .ZN(n731) );
  XNOR2_X1 U460 ( .A(n502), .B(n487), .ZN(n486) );
  INV_X1 U461 ( .A(G137), .ZN(n487) );
  INV_X1 U462 ( .A(KEYINPUT74), .ZN(n472) );
  XNOR2_X1 U463 ( .A(KEYINPUT17), .B(KEYINPUT78), .ZN(n503) );
  XNOR2_X1 U464 ( .A(n385), .B(n384), .ZN(n690) );
  INV_X1 U465 ( .A(KEYINPUT110), .ZN(n384) );
  INV_X1 U466 ( .A(KEYINPUT105), .ZN(n445) );
  INV_X1 U467 ( .A(KEYINPUT73), .ZN(n434) );
  NAND2_X1 U468 ( .A1(G214), .A2(n561), .ZN(n686) );
  NOR2_X1 U469 ( .A1(n558), .A2(n571), .ZN(n568) );
  XNOR2_X1 U470 ( .A(n521), .B(n439), .ZN(n640) );
  XNOR2_X1 U471 ( .A(n525), .B(n520), .ZN(n439) );
  NAND2_X1 U472 ( .A1(n485), .A2(n392), .ZN(n391) );
  INV_X1 U473 ( .A(G902), .ZN(n392) );
  NAND2_X1 U474 ( .A1(n559), .A2(G472), .ZN(n395) );
  XNOR2_X1 U475 ( .A(n402), .B(n596), .ZN(n401) );
  INV_X1 U476 ( .A(n666), .ZN(n440) );
  XNOR2_X1 U477 ( .A(n496), .B(KEYINPUT3), .ZN(n462) );
  XNOR2_X1 U478 ( .A(n389), .B(n388), .ZN(n387) );
  INV_X1 U479 ( .A(G113), .ZN(n496) );
  XNOR2_X1 U480 ( .A(n475), .B(n474), .ZN(n473) );
  XNOR2_X1 U481 ( .A(KEYINPUT24), .B(G140), .ZN(n475) );
  XNOR2_X1 U482 ( .A(G128), .B(G110), .ZN(n474) );
  XNOR2_X1 U483 ( .A(n546), .B(KEYINPUT76), .ZN(n476) );
  XNOR2_X1 U484 ( .A(G119), .B(G137), .ZN(n546) );
  XNOR2_X1 U485 ( .A(n544), .B(n545), .ZN(n548) );
  XNOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n545) );
  XNOR2_X1 U487 ( .A(KEYINPUT77), .B(G101), .ZN(n454) );
  INV_X1 U488 ( .A(KEYINPUT0), .ZN(n432) );
  NOR2_X2 U489 ( .A1(n367), .A2(n603), .ZN(n433) );
  INV_X1 U490 ( .A(KEYINPUT89), .ZN(n509) );
  XNOR2_X1 U491 ( .A(n566), .B(KEYINPUT103), .ZN(n582) );
  NAND2_X1 U492 ( .A1(n615), .A2(n400), .ZN(n572) );
  AND2_X1 U493 ( .A1(n493), .A2(G472), .ZN(n364) );
  XNOR2_X1 U494 ( .A(n460), .B(n366), .ZN(n728) );
  XNOR2_X1 U495 ( .A(n419), .B(n500), .ZN(n460) );
  XOR2_X1 U496 ( .A(G122), .B(KEYINPUT16), .Z(n500) );
  XNOR2_X1 U497 ( .A(n449), .B(n531), .ZN(n716) );
  XNOR2_X1 U498 ( .A(n450), .B(n535), .ZN(n449) );
  AND2_X1 U499 ( .A1(n684), .A2(n386), .ZN(n569) );
  INV_X1 U500 ( .A(n581), .ZN(n386) );
  XNOR2_X1 U501 ( .A(n478), .B(n477), .ZN(n745) );
  XNOR2_X1 U502 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n477) );
  INV_X1 U503 ( .A(n618), .ZN(n490) );
  XNOR2_X1 U504 ( .A(n610), .B(n464), .ZN(n463) );
  OR2_X1 U505 ( .A1(n612), .A2(n609), .ZN(n465) );
  INV_X1 U506 ( .A(KEYINPUT32), .ZN(n610) );
  INV_X1 U507 ( .A(n657), .ZN(n653) );
  NOR2_X1 U508 ( .A1(n396), .A2(n677), .ZN(n613) );
  XNOR2_X1 U509 ( .A(n625), .B(KEYINPUT107), .ZN(n744) );
  NAND2_X1 U510 ( .A1(n372), .A2(n369), .ZN(n368) );
  AND2_X1 U511 ( .A1(n375), .A2(n374), .ZN(n373) );
  AND2_X1 U512 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U513 ( .A(n713), .B(n712), .ZN(n714) );
  INV_X1 U514 ( .A(KEYINPUT56), .ZN(n479) );
  AND2_X1 U515 ( .A1(n376), .A2(n356), .ZN(n344) );
  XOR2_X1 U516 ( .A(n555), .B(n554), .Z(n345) );
  XOR2_X1 U517 ( .A(n501), .B(n502), .Z(n346) );
  INV_X1 U518 ( .A(n673), .ZN(n466) );
  XOR2_X1 U519 ( .A(n510), .B(n509), .Z(n347) );
  AND2_X1 U520 ( .A1(n677), .A2(n416), .ZN(n348) );
  AND2_X1 U521 ( .A1(n519), .A2(G210), .ZN(n349) );
  AND2_X1 U522 ( .A1(n440), .A2(n664), .ZN(n350) );
  INV_X1 U523 ( .A(G472), .ZN(n485) );
  XOR2_X1 U524 ( .A(n640), .B(n491), .Z(n351) );
  XOR2_X1 U525 ( .A(n616), .B(KEYINPUT108), .Z(n352) );
  AND2_X1 U526 ( .A1(n351), .A2(G475), .ZN(n353) );
  XOR2_X1 U527 ( .A(n559), .B(KEYINPUT62), .Z(n354) );
  XOR2_X1 U528 ( .A(n709), .B(n708), .Z(n355) );
  NOR2_X1 U529 ( .A1(G952), .A2(n704), .ZN(n721) );
  INV_X1 U530 ( .A(n721), .ZN(n382) );
  XOR2_X1 U531 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n356) );
  XOR2_X1 U532 ( .A(n637), .B(KEYINPUT85), .Z(n357) );
  INV_X1 U533 ( .A(G953), .ZN(n704) );
  NAND2_X1 U534 ( .A1(n358), .A2(n627), .ZN(n436) );
  NAND2_X1 U535 ( .A1(n684), .A2(n358), .ZN(n668) );
  NAND2_X1 U536 ( .A1(n695), .A2(n358), .ZN(n696) );
  XNOR2_X2 U537 ( .A(n483), .B(n352), .ZN(n358) );
  NAND2_X1 U538 ( .A1(n360), .A2(n425), .ZN(n423) );
  NAND2_X1 U539 ( .A1(n361), .A2(n424), .ZN(n360) );
  INV_X1 U540 ( .A(n426), .ZN(n361) );
  NAND2_X1 U541 ( .A1(n362), .A2(n494), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n363), .A2(n494), .ZN(n381) );
  NAND2_X1 U543 ( .A1(n364), .A2(n494), .ZN(n458) );
  NAND2_X1 U544 ( .A1(n365), .A2(G217), .ZN(n718) );
  NAND2_X1 U545 ( .A1(n365), .A2(G478), .ZN(n715) );
  NAND2_X1 U546 ( .A1(n365), .A2(G469), .ZN(n713) );
  XNOR2_X1 U547 ( .A(n366), .B(n497), .ZN(n498) );
  NOR2_X1 U548 ( .A1(n581), .A2(n367), .ZN(n654) );
  NAND2_X1 U549 ( .A1(n373), .A2(n368), .ZN(G60) );
  INV_X1 U550 ( .A(n356), .ZN(n370) );
  NAND2_X1 U551 ( .A1(n377), .A2(n376), .ZN(n371) );
  NAND2_X1 U552 ( .A1(n377), .A2(n344), .ZN(n374) );
  INV_X1 U553 ( .A(n588), .ZN(n590) );
  NAND2_X1 U554 ( .A1(n588), .A2(n686), .ZN(n428) );
  XNOR2_X2 U555 ( .A(n511), .B(n347), .ZN(n588) );
  NAND2_X1 U556 ( .A1(n383), .A2(n403), .ZN(n402) );
  XNOR2_X1 U557 ( .A(n458), .B(n354), .ZN(n457) );
  NAND2_X1 U558 ( .A1(n687), .A2(n686), .ZN(n385) );
  NAND2_X1 U559 ( .A1(n397), .A2(n466), .ZN(n558) );
  INV_X1 U560 ( .A(n397), .ZN(n396) );
  XNOR2_X1 U561 ( .A(n397), .B(KEYINPUT106), .ZN(n674) );
  XNOR2_X2 U562 ( .A(n467), .B(n345), .ZN(n397) );
  NAND2_X1 U563 ( .A1(n398), .A2(n677), .ZN(n682) );
  XNOR2_X2 U564 ( .A(n435), .B(n434), .ZN(n398) );
  XNOR2_X2 U565 ( .A(n731), .B(G146), .ZN(n399) );
  INV_X1 U566 ( .A(n417), .ZN(n400) );
  XNOR2_X2 U567 ( .A(n417), .B(KEYINPUT1), .ZN(n671) );
  XNOR2_X2 U568 ( .A(n513), .B(G469), .ZN(n417) );
  AND2_X1 U569 ( .A1(n430), .A2(n663), .ZN(n403) );
  AND2_X1 U570 ( .A1(n654), .A2(n406), .ZN(n405) );
  XNOR2_X1 U571 ( .A(n691), .B(KEYINPUT82), .ZN(n632) );
  NAND2_X1 U572 ( .A1(n409), .A2(n652), .ZN(n408) );
  NAND2_X1 U573 ( .A1(n583), .A2(KEYINPUT47), .ZN(n409) );
  NAND2_X1 U574 ( .A1(n412), .A2(n410), .ZN(n581) );
  INV_X1 U575 ( .A(n568), .ZN(n411) );
  AND2_X1 U576 ( .A1(n415), .A2(n413), .ZN(n412) );
  NOR2_X1 U577 ( .A1(n414), .A2(n417), .ZN(n413) );
  NOR2_X1 U578 ( .A1(n677), .A2(n416), .ZN(n414) );
  NAND2_X1 U579 ( .A1(n568), .A2(n348), .ZN(n415) );
  INV_X1 U580 ( .A(KEYINPUT28), .ZN(n416) );
  AND2_X2 U581 ( .A1(n470), .A2(n418), .ZN(n667) );
  INV_X1 U582 ( .A(n733), .ZN(n418) );
  NAND2_X1 U583 ( .A1(n470), .A2(n704), .ZN(n725) );
  XNOR2_X2 U584 ( .A(n429), .B(KEYINPUT45), .ZN(n470) );
  XNOR2_X1 U585 ( .A(n512), .B(n419), .ZN(n455) );
  NAND2_X1 U586 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U587 ( .A1(n744), .A2(KEYINPUT84), .ZN(n421) );
  NAND2_X1 U588 ( .A1(n426), .A2(KEYINPUT84), .ZN(n422) );
  AND2_X2 U589 ( .A1(n427), .A2(n636), .ZN(n494) );
  NAND2_X1 U590 ( .A1(n667), .A2(KEYINPUT2), .ZN(n427) );
  NAND2_X1 U591 ( .A1(n448), .A2(n459), .ZN(n429) );
  XNOR2_X1 U592 ( .A(n589), .B(KEYINPUT72), .ZN(n430) );
  XNOR2_X2 U593 ( .A(n433), .B(n432), .ZN(n630) );
  NOR2_X2 U594 ( .A1(n671), .A2(n670), .ZN(n435) );
  NOR2_X2 U595 ( .A1(G902), .A2(n711), .ZN(n513) );
  NAND2_X1 U596 ( .A1(n597), .A2(n653), .ZN(n478) );
  XNOR2_X1 U597 ( .A(n436), .B(n617), .ZN(n443) );
  NAND2_X1 U598 ( .A1(n443), .A2(n490), .ZN(n442) );
  NOR2_X1 U599 ( .A1(n653), .A2(n649), .ZN(n438) );
  OR2_X2 U600 ( .A1(n743), .A2(KEYINPUT44), .ZN(n619) );
  XNOR2_X1 U601 ( .A(n620), .B(KEYINPUT69), .ZN(n459) );
  NAND2_X1 U602 ( .A1(n743), .A2(KEYINPUT44), .ZN(n635) );
  XNOR2_X2 U603 ( .A(n442), .B(KEYINPUT35), .ZN(n743) );
  NAND2_X1 U604 ( .A1(n688), .A2(n466), .ZN(n446) );
  INV_X1 U605 ( .A(KEYINPUT19), .ZN(n447) );
  XNOR2_X1 U606 ( .A(n456), .B(n357), .ZN(G57) );
  NAND2_X1 U607 ( .A1(n457), .A2(n382), .ZN(n456) );
  NAND2_X1 U608 ( .A1(n471), .A2(n470), .ZN(n469) );
  XNOR2_X1 U609 ( .A(n733), .B(n472), .ZN(n471) );
  XNOR2_X1 U610 ( .A(n480), .B(n479), .ZN(G51) );
  NAND2_X1 U611 ( .A1(n481), .A2(n382), .ZN(n480) );
  XNOR2_X1 U612 ( .A(n482), .B(n355), .ZN(n481) );
  XNOR2_X2 U613 ( .A(n489), .B(G128), .ZN(n501) );
  XNOR2_X1 U614 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U615 ( .A(n639), .B(n638), .Z(n491) );
  XOR2_X1 U616 ( .A(n534), .B(n533), .Z(n492) );
  INV_X1 U617 ( .A(KEYINPUT103), .ZN(n565) );
  INV_X1 U618 ( .A(G478), .ZN(n537) );
  XNOR2_X1 U619 ( .A(n577), .B(KEYINPUT70), .ZN(n578) );
  XOR2_X1 U620 ( .A(KEYINPUT75), .B(n499), .Z(n519) );
  INV_X1 U621 ( .A(n552), .ZN(n636) );
  XNOR2_X1 U622 ( .A(n503), .B(n514), .ZN(n504) );
  XOR2_X1 U623 ( .A(KEYINPUT18), .B(n504), .Z(n506) );
  NAND2_X1 U624 ( .A1(G224), .A2(n704), .ZN(n505) );
  XNOR2_X1 U625 ( .A(n506), .B(n505), .ZN(n507) );
  AND2_X1 U626 ( .A1(G210), .A2(n561), .ZN(n510) );
  XOR2_X1 U627 ( .A(G131), .B(G140), .Z(n515) );
  NAND2_X1 U628 ( .A1(G227), .A2(n704), .ZN(n512) );
  INV_X1 U629 ( .A(n671), .ZN(n611) );
  XNOR2_X1 U630 ( .A(n544), .B(n515), .ZN(n732) );
  XNOR2_X1 U631 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U632 ( .A(n732), .B(n518), .Z(n521) );
  NAND2_X1 U633 ( .A1(G214), .A2(n519), .ZN(n520) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U635 ( .A(KEYINPUT98), .B(n524), .Z(n525) );
  NOR2_X1 U636 ( .A1(G902), .A2(n640), .ZN(n527) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  XNOR2_X1 U638 ( .A(n528), .B(KEYINPUT100), .ZN(n536) );
  INV_X1 U639 ( .A(n529), .ZN(n530) );
  XOR2_X1 U640 ( .A(n530), .B(KEYINPUT102), .Z(n531) );
  NAND2_X1 U641 ( .A1(G217), .A2(n549), .ZN(n535) );
  NAND2_X1 U642 ( .A1(G234), .A2(G237), .ZN(n539) );
  XNOR2_X1 U643 ( .A(n539), .B(KEYINPUT90), .ZN(n540) );
  XNOR2_X1 U644 ( .A(KEYINPUT14), .B(n540), .ZN(n541) );
  NAND2_X1 U645 ( .A1(G952), .A2(n541), .ZN(n701) );
  NOR2_X1 U646 ( .A1(G953), .A2(n701), .ZN(n601) );
  AND2_X1 U647 ( .A1(n541), .A2(G902), .ZN(n598) );
  NAND2_X1 U648 ( .A1(G953), .A2(n598), .ZN(n542) );
  NOR2_X1 U649 ( .A1(G900), .A2(n542), .ZN(n543) );
  NOR2_X1 U650 ( .A1(n601), .A2(n543), .ZN(n571) );
  XNOR2_X1 U651 ( .A(n548), .B(n547), .ZN(n551) );
  NAND2_X1 U652 ( .A1(n549), .A2(G221), .ZN(n550) );
  XNOR2_X1 U653 ( .A(n551), .B(n550), .ZN(n719) );
  NAND2_X1 U654 ( .A1(G234), .A2(n552), .ZN(n553) );
  XNOR2_X1 U655 ( .A(KEYINPUT20), .B(n553), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n556), .A2(G217), .ZN(n554) );
  NAND2_X1 U657 ( .A1(n556), .A2(G221), .ZN(n557) );
  XNOR2_X1 U658 ( .A(KEYINPUT21), .B(n557), .ZN(n673) );
  NAND2_X1 U659 ( .A1(n568), .A2(n622), .ZN(n560) );
  NOR2_X1 U660 ( .A1(n657), .A2(n560), .ZN(n562) );
  NAND2_X1 U661 ( .A1(n562), .A2(n686), .ZN(n591) );
  NOR2_X1 U662 ( .A1(n611), .A2(n591), .ZN(n563) );
  XNOR2_X1 U663 ( .A(n563), .B(KEYINPUT43), .ZN(n564) );
  NOR2_X1 U664 ( .A1(n588), .A2(n564), .ZN(n666) );
  XNOR2_X1 U665 ( .A(KEYINPUT38), .B(n590), .ZN(n687) );
  NOR2_X1 U666 ( .A1(n585), .A2(n584), .ZN(n688) );
  NAND2_X1 U667 ( .A1(n690), .A2(n688), .ZN(n567) );
  XNOR2_X1 U668 ( .A(KEYINPUT42), .B(n569), .ZN(n746) );
  INV_X1 U669 ( .A(n687), .ZN(n576) );
  NAND2_X1 U670 ( .A1(n677), .A2(n686), .ZN(n570) );
  XOR2_X1 U671 ( .A(n570), .B(KEYINPUT30), .Z(n575) );
  INV_X1 U672 ( .A(n571), .ZN(n573) );
  XNOR2_X1 U673 ( .A(KEYINPUT95), .B(n572), .ZN(n626) );
  AND2_X1 U674 ( .A1(n573), .A2(n626), .ZN(n574) );
  NAND2_X1 U675 ( .A1(n575), .A2(n574), .ZN(n586) );
  XNOR2_X1 U676 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n577) );
  NOR2_X1 U677 ( .A1(n746), .A2(n745), .ZN(n580) );
  NOR2_X1 U678 ( .A1(n584), .A2(n582), .ZN(n649) );
  NAND2_X1 U679 ( .A1(n654), .A2(n691), .ZN(n583) );
  NAND2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n618) );
  NOR2_X1 U681 ( .A1(n586), .A2(n618), .ZN(n587) );
  NAND2_X1 U682 ( .A1(n588), .A2(n587), .ZN(n652) );
  OR2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U684 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n592) );
  XNOR2_X1 U685 ( .A(n593), .B(n592), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n594), .A2(n611), .ZN(n663) );
  NAND2_X1 U687 ( .A1(n649), .A2(n597), .ZN(n664) );
  NOR2_X1 U688 ( .A1(G898), .A2(n704), .ZN(n727) );
  NAND2_X1 U689 ( .A1(n598), .A2(n727), .ZN(n599) );
  XNOR2_X1 U690 ( .A(KEYINPUT91), .B(n599), .ZN(n600) );
  NOR2_X1 U691 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U692 ( .A(n602), .B(KEYINPUT92), .ZN(n603) );
  XNOR2_X1 U693 ( .A(KEYINPUT22), .B(KEYINPUT65), .ZN(n604) );
  INV_X1 U694 ( .A(n622), .ZN(n606) );
  NAND2_X1 U695 ( .A1(n674), .A2(n606), .ZN(n607) );
  NOR2_X1 U696 ( .A1(n671), .A2(n607), .ZN(n608) );
  XOR2_X1 U697 ( .A(KEYINPUT80), .B(n608), .Z(n609) );
  NAND2_X1 U698 ( .A1(n613), .A2(n624), .ZN(n647) );
  XOR2_X1 U699 ( .A(KEYINPUT34), .B(KEYINPUT79), .Z(n614) );
  XNOR2_X1 U700 ( .A(KEYINPUT71), .B(n614), .ZN(n617) );
  INV_X1 U701 ( .A(n630), .ZN(n627) );
  INV_X1 U702 ( .A(n615), .ZN(n670) );
  XNOR2_X1 U703 ( .A(KEYINPUT33), .B(KEYINPUT87), .ZN(n616) );
  NOR2_X2 U704 ( .A1(n621), .A2(n619), .ZN(n620) );
  NOR2_X1 U705 ( .A1(n622), .A2(n674), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  AND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n629) );
  INV_X1 U708 ( .A(n677), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n642) );
  NOR2_X1 U710 ( .A1(n682), .A2(n630), .ZN(n631) );
  XNOR2_X1 U711 ( .A(n631), .B(KEYINPUT31), .ZN(n659) );
  NAND2_X1 U712 ( .A1(n642), .A2(n659), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT66), .B(KEYINPUT123), .Z(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT122), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n657), .A2(n642), .ZN(n641) );
  XOR2_X1 U718 ( .A(G104), .B(n641), .Z(G6) );
  INV_X1 U719 ( .A(n649), .ZN(n660) );
  NOR2_X1 U720 ( .A1(n642), .A2(n660), .ZN(n646) );
  XOR2_X1 U721 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n644) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT27), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(G9) );
  XNOR2_X1 U725 ( .A(G110), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n648), .B(n647), .ZN(G12) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U728 ( .A1(n649), .A2(n654), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(G30) );
  XNOR2_X1 U730 ( .A(G143), .B(n652), .ZN(G45) );
  XOR2_X1 U731 ( .A(G146), .B(KEYINPUT115), .Z(n656) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(G48) );
  NOR2_X1 U734 ( .A1(n657), .A2(n659), .ZN(n658) );
  XOR2_X1 U735 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U737 ( .A(G116), .B(n661), .Z(G18) );
  XOR2_X1 U738 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(KEYINPUT116), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(n664), .ZN(G36) );
  XOR2_X1 U742 ( .A(G140), .B(n666), .Z(G42) );
  XNOR2_X1 U743 ( .A(KEYINPUT2), .B(n667), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT50), .B(n672), .ZN(n680) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n676) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U752 ( .A(KEYINPUT51), .B(n683), .Z(n685) );
  NAND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n697) );
  OR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U758 ( .A(n694), .B(KEYINPUT118), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U760 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(KEYINPUT119), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n702), .B(KEYINPUT120), .ZN(n703) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT121), .ZN(n706) );
  XNOR2_X1 U765 ( .A(KEYINPUT53), .B(n706), .ZN(G75) );
  XOR2_X1 U766 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n709) );
  XNOR2_X1 U767 ( .A(n707), .B(KEYINPUT86), .ZN(n708) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n710) );
  NOR2_X1 U769 ( .A1(n721), .A2(n714), .ZN(G54) );
  XNOR2_X1 U770 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n721), .A2(n717), .ZN(G63) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(G66) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n722) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n722), .ZN(n723) );
  NAND2_X1 U776 ( .A1(n723), .A2(G898), .ZN(n724) );
  NAND2_X1 U777 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U778 ( .A(n726), .B(KEYINPUT125), .ZN(n730) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U780 ( .A(n730), .B(n729), .Z(G69) );
  XOR2_X1 U781 ( .A(n731), .B(n732), .Z(n736) );
  XOR2_X1 U782 ( .A(n733), .B(n736), .Z(n734) );
  XNOR2_X1 U783 ( .A(KEYINPUT126), .B(n734), .ZN(n735) );
  NOR2_X1 U784 ( .A1(G953), .A2(n735), .ZN(n740) );
  XNOR2_X1 U785 ( .A(G227), .B(n736), .ZN(n738) );
  NAND2_X1 U786 ( .A1(G900), .A2(G953), .ZN(n737) );
  NOR2_X1 U787 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U788 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n741), .Z(G72) );
  XNOR2_X1 U790 ( .A(G119), .B(n742), .ZN(G21) );
  XOR2_X1 U791 ( .A(n743), .B(G122), .Z(G24) );
  XOR2_X1 U792 ( .A(n744), .B(G101), .Z(G3) );
  XOR2_X1 U793 ( .A(n745), .B(G131), .Z(G33) );
  XOR2_X1 U794 ( .A(G137), .B(n746), .Z(G39) );
endmodule

