

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(G164), .A2(G1384), .ZN(n720) );
  INV_X1 U557 ( .A(n645), .ZN(n652) );
  AND2_X1 U558 ( .A1(n931), .A2(n744), .ZN(n522) );
  OR2_X1 U559 ( .A1(n732), .A2(n522), .ZN(n523) );
  XNOR2_X1 U560 ( .A(n594), .B(KEYINPUT26), .ZN(n604) );
  NOR2_X2 U561 ( .A1(n593), .A2(n719), .ZN(n645) );
  INV_X1 U562 ( .A(KEYINPUT103), .ZN(n693) );
  OR2_X1 U563 ( .A1(n733), .A2(n523), .ZN(n747) );
  NOR2_X1 U564 ( .A1(G651), .A2(n571), .ZN(n772) );
  NOR2_X1 U565 ( .A1(n603), .A2(n602), .ZN(n918) );
  INV_X1 U566 ( .A(G2104), .ZN(n527) );
  NOR2_X2 U567 ( .A1(G2105), .A2(n527), .ZN(n888) );
  NAND2_X1 U568 ( .A1(G102), .A2(n888), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n524), .Z(n889) );
  NAND2_X1 U571 ( .A1(G138), .A2(n889), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U573 ( .A1(n527), .A2(G2105), .ZN(n528) );
  XNOR2_X1 U574 ( .A(n528), .B(KEYINPUT65), .ZN(n892) );
  NAND2_X1 U575 ( .A1(n892), .A2(G126), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U577 ( .A(KEYINPUT66), .B(n529), .Z(n893) );
  NAND2_X1 U578 ( .A1(G114), .A2(n893), .ZN(n530) );
  NAND2_X1 U579 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U580 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U581 ( .A1(n893), .A2(G113), .ZN(n534) );
  XOR2_X1 U582 ( .A(n534), .B(KEYINPUT67), .Z(n537) );
  NAND2_X1 U583 ( .A1(G101), .A2(n888), .ZN(n535) );
  XOR2_X1 U584 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U586 ( .A1(G137), .A2(n889), .ZN(n539) );
  NAND2_X1 U587 ( .A1(G125), .A2(n892), .ZN(n538) );
  NAND2_X1 U588 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X2 U589 ( .A1(n541), .A2(n540), .ZN(G160) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n571) );
  NAND2_X1 U591 ( .A1(G52), .A2(n772), .ZN(n544) );
  INV_X1 U592 ( .A(G651), .ZN(n545) );
  NOR2_X1 U593 ( .A1(G543), .A2(n545), .ZN(n542) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n542), .Z(n778) );
  NAND2_X1 U595 ( .A1(G64), .A2(n778), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n551) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n777) );
  NAND2_X1 U598 ( .A1(G90), .A2(n777), .ZN(n547) );
  NOR2_X1 U599 ( .A1(n571), .A2(n545), .ZN(n774) );
  NAND2_X1 U600 ( .A1(G77), .A2(n774), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT68), .B(n548), .Z(n549) );
  XNOR2_X1 U603 ( .A(KEYINPUT9), .B(n549), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(G171) );
  INV_X1 U605 ( .A(G171), .ZN(G301) );
  NAND2_X1 U606 ( .A1(G89), .A2(n777), .ZN(n552) );
  XOR2_X1 U607 ( .A(KEYINPUT4), .B(n552), .Z(n553) );
  XNOR2_X1 U608 ( .A(n553), .B(KEYINPUT75), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G76), .A2(n774), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G51), .A2(n772), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G63), .A2(n778), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U617 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G88), .A2(n777), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G75), .A2(n774), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n778), .A2(G62), .ZN(n565) );
  XOR2_X1 U623 ( .A(KEYINPUT84), .B(n565), .Z(n566) );
  NOR2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n772), .A2(G50), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(G303) );
  INV_X1 U627 ( .A(G303), .ZN(G166) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n570) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT80), .ZN(n576) );
  NAND2_X1 U630 ( .A1(G49), .A2(n772), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G87), .A2(n571), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n778), .A2(n574), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U635 ( .A(KEYINPUT81), .B(n577), .Z(G288) );
  NAND2_X1 U636 ( .A1(G73), .A2(n774), .ZN(n578) );
  XNOR2_X1 U637 ( .A(n578), .B(KEYINPUT2), .ZN(n586) );
  NAND2_X1 U638 ( .A1(n777), .A2(G86), .ZN(n579) );
  XNOR2_X1 U639 ( .A(n579), .B(KEYINPUT82), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G61), .A2(n778), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U642 ( .A1(G48), .A2(n772), .ZN(n582) );
  XNOR2_X1 U643 ( .A(KEYINPUT83), .B(n582), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U646 ( .A1(G85), .A2(n777), .ZN(n588) );
  NAND2_X1 U647 ( .A1(G72), .A2(n774), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U649 ( .A1(G47), .A2(n772), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G60), .A2(n778), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U652 ( .A1(n592), .A2(n591), .ZN(G290) );
  INV_X1 U653 ( .A(KEYINPUT29), .ZN(n644) );
  INV_X1 U654 ( .A(n720), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n719) );
  NAND2_X1 U656 ( .A1(n645), .A2(G1996), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n777), .A2(G81), .ZN(n595) );
  XNOR2_X1 U658 ( .A(n595), .B(KEYINPUT12), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G68), .A2(n774), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U661 ( .A(n598), .B(KEYINPUT13), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G43), .A2(n772), .ZN(n599) );
  NAND2_X1 U663 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U664 ( .A1(n778), .A2(G56), .ZN(n601) );
  XOR2_X1 U665 ( .A(KEYINPUT14), .B(n601), .Z(n602) );
  NAND2_X1 U666 ( .A1(n604), .A2(n918), .ZN(n607) );
  NAND2_X1 U667 ( .A1(G1341), .A2(n652), .ZN(n605) );
  XNOR2_X1 U668 ( .A(n605), .B(KEYINPUT97), .ZN(n606) );
  NOR2_X1 U669 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U670 ( .A(KEYINPUT64), .ZN(n608) );
  XNOR2_X1 U671 ( .A(n609), .B(n608), .ZN(n624) );
  NAND2_X1 U672 ( .A1(G79), .A2(n774), .ZN(n610) );
  XNOR2_X1 U673 ( .A(n610), .B(KEYINPUT74), .ZN(n617) );
  NAND2_X1 U674 ( .A1(G54), .A2(n772), .ZN(n612) );
  NAND2_X1 U675 ( .A1(G66), .A2(n778), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U677 ( .A1(G92), .A2(n777), .ZN(n613) );
  XNOR2_X1 U678 ( .A(KEYINPUT73), .B(n613), .ZN(n614) );
  NOR2_X1 U679 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U680 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U681 ( .A(KEYINPUT15), .B(n618), .Z(n923) );
  OR2_X1 U682 ( .A1(n624), .A2(n923), .ZN(n623) );
  AND2_X1 U683 ( .A1(n645), .A2(G2067), .ZN(n619) );
  XOR2_X1 U684 ( .A(n619), .B(KEYINPUT98), .Z(n621) );
  NAND2_X1 U685 ( .A1(n652), .A2(G1348), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U687 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U688 ( .A1(n624), .A2(n923), .ZN(n625) );
  NAND2_X1 U689 ( .A1(n626), .A2(n625), .ZN(n638) );
  NAND2_X1 U690 ( .A1(G53), .A2(n772), .ZN(n628) );
  NAND2_X1 U691 ( .A1(G65), .A2(n778), .ZN(n627) );
  NAND2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U693 ( .A1(G91), .A2(n777), .ZN(n630) );
  NAND2_X1 U694 ( .A1(G78), .A2(n774), .ZN(n629) );
  NAND2_X1 U695 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U696 ( .A1(n632), .A2(n631), .ZN(n927) );
  NAND2_X1 U697 ( .A1(G2072), .A2(n645), .ZN(n633) );
  XNOR2_X1 U698 ( .A(n633), .B(KEYINPUT96), .ZN(n634) );
  XNOR2_X1 U699 ( .A(KEYINPUT27), .B(n634), .ZN(n636) );
  INV_X1 U700 ( .A(G1956), .ZN(n836) );
  NOR2_X1 U701 ( .A1(n645), .A2(n836), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U703 ( .A1(n927), .A2(n639), .ZN(n637) );
  NAND2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U705 ( .A1(n927), .A2(n639), .ZN(n640) );
  XOR2_X1 U706 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  AND2_X1 U707 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n644), .B(n643), .ZN(n650) );
  NAND2_X1 U709 ( .A1(G1961), .A2(n652), .ZN(n647) );
  XOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NAND2_X1 U711 ( .A1(n645), .A2(n948), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n657) );
  NOR2_X1 U713 ( .A1(G301), .A2(n657), .ZN(n648) );
  XOR2_X1 U714 ( .A(KEYINPUT95), .B(n648), .Z(n649) );
  NOR2_X2 U715 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U716 ( .A(n651), .B(KEYINPUT99), .ZN(n662) );
  NAND2_X1 U717 ( .A1(G8), .A2(n652), .ZN(n698) );
  NOR2_X1 U718 ( .A1(G1966), .A2(n698), .ZN(n675) );
  NOR2_X1 U719 ( .A1(G2084), .A2(n652), .ZN(n672) );
  NOR2_X1 U720 ( .A1(n675), .A2(n672), .ZN(n653) );
  NAND2_X1 U721 ( .A1(G8), .A2(n653), .ZN(n654) );
  XNOR2_X1 U722 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U723 ( .A1(G168), .A2(n655), .ZN(n656) );
  XOR2_X1 U724 ( .A(KEYINPUT100), .B(n656), .Z(n659) );
  NAND2_X1 U725 ( .A1(G301), .A2(n657), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(KEYINPUT31), .B(n660), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n673) );
  NAND2_X1 U729 ( .A1(n673), .A2(G286), .ZN(n670) );
  INV_X1 U730 ( .A(G8), .ZN(n668) );
  NOR2_X1 U731 ( .A1(G1971), .A2(n698), .ZN(n663) );
  XNOR2_X1 U732 ( .A(KEYINPUT101), .B(n663), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n652), .ZN(n664) );
  NOR2_X1 U734 ( .A1(G166), .A2(n664), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  OR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(n671), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U739 ( .A1(G8), .A2(n672), .ZN(n677) );
  INV_X1 U740 ( .A(n673), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n692) );
  NOR2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n934) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n929) );
  NOR2_X1 U746 ( .A1(n934), .A2(n929), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n692), .A2(n680), .ZN(n683) );
  INV_X1 U748 ( .A(n698), .ZN(n681) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n935) );
  AND2_X1 U750 ( .A1(n681), .A2(n935), .ZN(n682) );
  AND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(KEYINPUT33), .A2(n684), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n934), .A2(KEYINPUT33), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n685), .A2(n698), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n915) );
  AND2_X1 U757 ( .A1(n688), .A2(n915), .ZN(n702) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U759 ( .A1(G8), .A2(n689), .ZN(n690) );
  XNOR2_X1 U760 ( .A(n690), .B(KEYINPUT102), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n695), .A2(n698), .ZN(n700) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n696) );
  XOR2_X1 U765 ( .A(n696), .B(KEYINPUT24), .Z(n697) );
  OR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n733) );
  NAND2_X1 U769 ( .A1(G95), .A2(n888), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G131), .A2(n889), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n892), .A2(G119), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G107), .A2(n893), .ZN(n705) );
  NAND2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n883) );
  INV_X1 U776 ( .A(G1991), .ZN(n954) );
  NOR2_X1 U777 ( .A1(n883), .A2(n954), .ZN(n718) );
  NAND2_X1 U778 ( .A1(G129), .A2(n892), .ZN(n709) );
  XNOR2_X1 U779 ( .A(n709), .B(KEYINPUT92), .ZN(n716) );
  NAND2_X1 U780 ( .A1(G141), .A2(n889), .ZN(n711) );
  NAND2_X1 U781 ( .A1(G117), .A2(n893), .ZN(n710) );
  NAND2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n888), .A2(G105), .ZN(n712) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U785 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U786 ( .A1(n716), .A2(n715), .ZN(n901) );
  AND2_X1 U787 ( .A1(n901), .A2(G1996), .ZN(n717) );
  OR2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n971) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n744) );
  AND2_X1 U790 ( .A1(n971), .A2(n744), .ZN(n736) );
  XNOR2_X1 U791 ( .A(KEYINPUT93), .B(n736), .ZN(n730) );
  XNOR2_X1 U792 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NAND2_X1 U793 ( .A1(G104), .A2(n888), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G140), .A2(n889), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n723), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n892), .A2(G128), .ZN(n725) );
  NAND2_X1 U798 ( .A1(G116), .A2(n893), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U800 ( .A(KEYINPUT35), .B(n726), .Z(n727) );
  NOR2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n729), .ZN(n905) );
  NOR2_X1 U803 ( .A1(n742), .A2(n905), .ZN(n970) );
  NAND2_X1 U804 ( .A1(n744), .A2(n970), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n730), .A2(n740), .ZN(n731) );
  XNOR2_X1 U806 ( .A(n731), .B(KEYINPUT94), .ZN(n732) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n931) );
  AND2_X1 U808 ( .A1(n954), .A2(n883), .ZN(n984) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n984), .A2(n734), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U812 ( .A1(G1996), .A2(n901), .ZN(n977) );
  NOR2_X1 U813 ( .A1(n737), .A2(n977), .ZN(n738) );
  XNOR2_X1 U814 ( .A(n738), .B(KEYINPUT104), .ZN(n739) );
  XNOR2_X1 U815 ( .A(n739), .B(KEYINPUT39), .ZN(n741) );
  NAND2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n742), .A2(n905), .ZN(n979) );
  NAND2_X1 U818 ( .A1(n743), .A2(n979), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U821 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U822 ( .A1(G111), .A2(n893), .ZN(n755) );
  NAND2_X1 U823 ( .A1(G99), .A2(n888), .ZN(n750) );
  NAND2_X1 U824 ( .A1(G135), .A2(n889), .ZN(n749) );
  NAND2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n892), .A2(G123), .ZN(n751) );
  XOR2_X1 U827 ( .A(KEYINPUT18), .B(n751), .Z(n752) );
  NOR2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U830 ( .A(KEYINPUT77), .B(n756), .Z(n981) );
  XNOR2_X1 U831 ( .A(G2096), .B(n981), .ZN(n757) );
  OR2_X1 U832 ( .A1(G2100), .A2(n757), .ZN(G156) );
  INV_X1 U833 ( .A(G132), .ZN(G219) );
  INV_X1 U834 ( .A(G96), .ZN(G221) );
  INV_X1 U835 ( .A(G57), .ZN(G237) );
  NAND2_X1 U836 ( .A1(G94), .A2(G452), .ZN(n758) );
  XNOR2_X1 U837 ( .A(n758), .B(KEYINPUT69), .ZN(G173) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n761) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n759) );
  XOR2_X1 U840 ( .A(n759), .B(KEYINPUT10), .Z(n818) );
  NAND2_X1 U841 ( .A1(G567), .A2(n818), .ZN(n760) );
  XNOR2_X1 U842 ( .A(n761), .B(n760), .ZN(G234) );
  NAND2_X1 U843 ( .A1(n918), .A2(G860), .ZN(G153) );
  NAND2_X1 U844 ( .A1(G868), .A2(G301), .ZN(n763) );
  INV_X1 U845 ( .A(G868), .ZN(n797) );
  NAND2_X1 U846 ( .A1(n923), .A2(n797), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n763), .A2(n762), .ZN(G284) );
  XOR2_X1 U848 ( .A(n927), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U849 ( .A1(G299), .A2(G868), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G286), .A2(n797), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(G297) );
  INV_X1 U852 ( .A(G860), .ZN(n785) );
  NAND2_X1 U853 ( .A1(n785), .A2(G559), .ZN(n766) );
  INV_X1 U854 ( .A(n923), .ZN(n783) );
  NAND2_X1 U855 ( .A1(n766), .A2(n783), .ZN(n767) );
  XNOR2_X1 U856 ( .A(n767), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(n923), .A2(n797), .ZN(n768) );
  XOR2_X1 U858 ( .A(KEYINPUT76), .B(n768), .Z(n769) );
  NOR2_X1 U859 ( .A1(G559), .A2(n769), .ZN(n771) );
  AND2_X1 U860 ( .A1(n797), .A2(n918), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(G282) );
  NAND2_X1 U862 ( .A1(G55), .A2(n772), .ZN(n773) );
  XNOR2_X1 U863 ( .A(n773), .B(KEYINPUT78), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n774), .A2(G80), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G93), .A2(n777), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G67), .A2(n778), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n796) );
  NAND2_X1 U870 ( .A1(G559), .A2(n783), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(n918), .ZN(n794) );
  NAND2_X1 U872 ( .A1(n785), .A2(n794), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT79), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n796), .B(n787), .ZN(G145) );
  XOR2_X1 U875 ( .A(G303), .B(n796), .Z(n793) );
  XNOR2_X1 U876 ( .A(G299), .B(G305), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n788), .B(G288), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT85), .B(n789), .ZN(n791) );
  XNOR2_X1 U879 ( .A(G290), .B(KEYINPUT19), .ZN(n790) );
  XNOR2_X1 U880 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n793), .B(n792), .ZN(n858) );
  XOR2_X1 U882 ( .A(n858), .B(n794), .Z(n795) );
  NOR2_X1 U883 ( .A1(n797), .A2(n795), .ZN(n799) );
  AND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(G295) );
  NAND2_X1 U886 ( .A1(G2078), .A2(G2084), .ZN(n800) );
  XOR2_X1 U887 ( .A(KEYINPUT20), .B(n800), .Z(n801) );
  NAND2_X1 U888 ( .A1(n801), .A2(G2090), .ZN(n802) );
  XNOR2_X1 U889 ( .A(n802), .B(KEYINPUT21), .ZN(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT86), .B(n803), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G2072), .A2(n804), .ZN(G158) );
  XOR2_X1 U892 ( .A(KEYINPUT87), .B(G44), .Z(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT3), .B(n805), .ZN(G218) );
  XNOR2_X1 U894 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U895 ( .A1(G69), .A2(G120), .ZN(n806) );
  NOR2_X1 U896 ( .A1(G237), .A2(n806), .ZN(n807) );
  NAND2_X1 U897 ( .A1(G108), .A2(n807), .ZN(n823) );
  NAND2_X1 U898 ( .A1(n823), .A2(G567), .ZN(n815) );
  NOR2_X1 U899 ( .A1(G219), .A2(G220), .ZN(n808) );
  XOR2_X1 U900 ( .A(KEYINPUT88), .B(n808), .Z(n809) );
  XNOR2_X1 U901 ( .A(n809), .B(KEYINPUT22), .ZN(n810) );
  NOR2_X1 U902 ( .A1(G218), .A2(n810), .ZN(n811) );
  XNOR2_X1 U903 ( .A(n811), .B(KEYINPUT89), .ZN(n812) );
  NOR2_X1 U904 ( .A1(G221), .A2(n812), .ZN(n813) );
  XOR2_X1 U905 ( .A(KEYINPUT90), .B(n813), .Z(n824) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n824), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n825) );
  NAND2_X1 U908 ( .A1(G483), .A2(G661), .ZN(n816) );
  NOR2_X1 U909 ( .A1(n825), .A2(n816), .ZN(n820) );
  NAND2_X1 U910 ( .A1(n820), .A2(G36), .ZN(n817) );
  XOR2_X1 U911 ( .A(KEYINPUT91), .B(n817), .Z(G176) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n818), .ZN(G217) );
  INV_X1 U913 ( .A(n818), .ZN(G223) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U915 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n822), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n825), .ZN(G319) );
  XNOR2_X1 U925 ( .A(G1348), .B(G2454), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n826), .B(G2430), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n827), .B(G1341), .ZN(n833) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n829) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n831) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n834), .A2(G14), .ZN(n835) );
  XNOR2_X1 U935 ( .A(KEYINPUT105), .B(n835), .ZN(G401) );
  XNOR2_X1 U936 ( .A(G1961), .B(G2474), .ZN(n846) );
  XOR2_X1 U937 ( .A(G1976), .B(G1981), .Z(n838) );
  XOR2_X1 U938 ( .A(G1966), .B(n836), .Z(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U940 ( .A(G1971), .B(G1986), .Z(n840) );
  XOR2_X1 U941 ( .A(G1996), .B(n954), .Z(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U943 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(G229) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2090), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n847), .B(KEYINPUT107), .ZN(n857) );
  XOR2_X1 U949 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2678), .B(G2096), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U952 ( .A(G2100), .B(G2078), .Z(n851) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U954 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U955 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT43), .B(KEYINPUT42), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U959 ( .A(n923), .B(n918), .Z(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n860) );
  XOR2_X1 U961 ( .A(G301), .B(n858), .Z(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(G286), .ZN(n864) );
  NOR2_X1 U965 ( .A1(G37), .A2(n864), .ZN(G397) );
  NAND2_X1 U966 ( .A1(G100), .A2(n888), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G136), .A2(n889), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G124), .A2(n892), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U971 ( .A1(G112), .A2(n893), .ZN(n868) );
  NAND2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G106), .A2(n888), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G142), .A2(n889), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT45), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G130), .A2(n892), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G118), .A2(n893), .ZN(n877) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n877), .ZN(n878) );
  NOR2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n887) );
  XOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U984 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n880) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(n882), .B(KEYINPUT113), .Z(n885) );
  XNOR2_X1 U987 ( .A(n883), .B(KEYINPUT112), .ZN(n884) );
  XNOR2_X1 U988 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n900) );
  NAND2_X1 U990 ( .A1(G103), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U993 ( .A1(n892), .A2(G127), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G115), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n972) );
  XNOR2_X1 U998 ( .A(n981), .B(n972), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(G162), .B(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(G164), .B(G160), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT116), .B(n909), .ZN(G395) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n911), .ZN(n912) );
  AND2_X1 U1010 ( .A1(G319), .A2(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(G16), .B(KEYINPUT56), .ZN(n943) );
  XNOR2_X1 U1016 ( .A(G1966), .B(G168), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT57), .ZN(n922) );
  XOR2_X1 U1019 ( .A(n918), .B(G1341), .Z(n920) );
  XOR2_X1 U1020 ( .A(G171), .B(G1961), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(G1348), .B(n923), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT122), .B(n924), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n941) );
  XOR2_X1 U1026 ( .A(n927), .B(G1956), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n933) );
  AND2_X1 U1028 ( .A1(G303), .A2(G1971), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(KEYINPUT123), .B(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(n939), .B(KEYINPUT124), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(n944), .B(KEYINPUT125), .ZN(n969) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G32), .B(G1996), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G27), .B(n948), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1047 ( .A(G25), .B(n954), .Z(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(n958), .B(KEYINPUT121), .ZN(n963) );
  XNOR2_X1 U1051 ( .A(G2084), .B(G34), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n959), .B(KEYINPUT54), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT55), .B(n964), .Z(n966) );
  INV_X1 U1057 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n967), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n997) );
  OR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n991) );
  XOR2_X1 U1062 ( .A(G2072), .B(n972), .Z(n974) );
  XOR2_X1 U1063 ( .A(G164), .B(G2078), .Z(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(KEYINPUT50), .B(n975), .ZN(n989) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(KEYINPUT51), .B(n978), .Z(n980) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n987) );
  XNOR2_X1 U1070 ( .A(G160), .B(G2084), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(KEYINPUT119), .B(n985), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n992), .ZN(n994) );
  INV_X1 U1078 ( .A(KEYINPUT55), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n995), .A2(G29), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(n997), .A2(n996), .ZN(n1022) );
  XOR2_X1 U1082 ( .A(G1976), .B(G23), .Z(n999) );
  XOR2_X1 U1083 ( .A(G1971), .B(G22), .Z(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G24), .B(G1986), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1087 ( .A(KEYINPUT58), .B(n1002), .Z(n1018) );
  XOR2_X1 U1088 ( .A(G1961), .B(G5), .Z(n1013) );
  XOR2_X1 U1089 ( .A(G4), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1004), .B(n1003), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(G20), .B(G1956), .Z(n1008) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G6), .B(G1981), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1011), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(G16), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

