//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  AOI21_X1  g002(.A(G8gat), .B1(new_n203), .B2(KEYINPUT90), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n206), .C1(KEYINPUT90), .C2(G8gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT17), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  OR2_X1    g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT88), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT89), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n213), .A2(new_n212), .A3(new_n214), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n215), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n215), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n211), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n229), .B(new_n211), .C1(new_n231), .C2(new_n225), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n210), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n229), .B1(new_n231), .B2(new_n225), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(new_n209), .A3(new_n208), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n237), .ZN(new_n241));
  INV_X1    g040(.A(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n210), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n237), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n235), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248));
  XOR2_X1   g047(.A(G169gat), .B(G197gat), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n254), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n256), .A3(new_n250), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n248), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n261), .A2(KEYINPUT12), .A3(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n247), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n260), .A2(new_n262), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n240), .A2(new_n264), .A3(new_n241), .A4(new_n246), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(G169gat), .A2(G176gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(KEYINPUT23), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT64), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  MUX2_X1   g071(.A(KEYINPUT24), .B(new_n271), .S(new_n272), .Z(new_n273));
  INV_X1    g072(.A(G169gat), .ZN(new_n274));
  INV_X1    g073(.A(G176gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(KEYINPUT23), .B2(new_n268), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT27), .B(G183gat), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n268), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(KEYINPUT26), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n276), .B2(KEYINPUT26), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n290), .A2(new_n291), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT25), .B1(new_n273), .B2(new_n279), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(new_n273), .A3(new_n270), .A4(new_n277), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n283), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n299));
  INV_X1    g098(.A(G127gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G134gat), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n300), .A2(G134gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(KEYINPUT66), .B(G134gat), .Z(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n304), .A2(G127gat), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n297), .A2(KEYINPUT1), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT69), .B1(new_n296), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n310), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n316), .B(KEYINPUT34), .Z(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n315), .ZN(new_n318));
  INV_X1    g117(.A(new_n314), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT33), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G15gat), .B(G43gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT70), .ZN(new_n325));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n320), .B(KEYINPUT32), .C1(new_n322), .C2(new_n327), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n317), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n329), .A3(KEYINPUT72), .A4(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G141gat), .B(G148gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT22), .ZN(new_n350));
  XNOR2_X1  g149(.A(G211gat), .B(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  INV_X1    g153(.A(G218gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n351), .B(new_n349), .C1(KEYINPUT22), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT73), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n345), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT84), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(new_n362), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n353), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT3), .B1(new_n365), .B2(new_n347), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n360), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G228gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT3), .B1(new_n358), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n361), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n375), .A2(G228gat), .A3(G233gat), .A4(new_n360), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G22gat), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n370), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(G78gat), .B(G106gat), .Z(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT82), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT31), .B(G50gat), .Z(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n381), .A2(KEYINPUT83), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n381), .B2(KEYINPUT83), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n329), .A2(new_n330), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n316), .B(KEYINPUT34), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n335), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n359), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n296), .A2(new_n371), .ZN(new_n395));
  INV_X1    g194(.A(G226gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n369), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n369), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n296), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(KEYINPUT75), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n394), .B(new_n397), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n296), .A2(new_n347), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n399), .B1(new_n403), .B2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n359), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G8gat), .B(G36gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT76), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  INV_X1    g212(.A(new_n411), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n406), .A2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n310), .A2(new_n345), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(KEYINPUT78), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n310), .A2(new_n345), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n420), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n421), .A2(new_n418), .A3(KEYINPUT4), .A4(new_n424), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n310), .B(KEYINPUT77), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n346), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G225gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT77), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n310), .B(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n421), .B(new_n424), .C1(new_n438), .C2(new_n361), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n434), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n422), .B2(KEYINPUT4), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n432), .B(new_n442), .C1(new_n425), .C2(KEYINPUT4), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT79), .B1(new_n440), .B2(KEYINPUT5), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n436), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(G1gat), .B(G29gat), .Z(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n449), .B(new_n450), .Z(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453));
  INV_X1    g252(.A(new_n451), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n436), .B(new_n454), .C1(new_n444), .C2(new_n445), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n417), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n393), .A2(new_n459), .A3(KEYINPUT35), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n391), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n390), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n335), .A3(new_n463), .A4(new_n389), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT35), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n335), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n335), .A2(new_n392), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(KEYINPUT36), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n457), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n411), .B1(new_n407), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n474), .B2(new_n407), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT38), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n404), .B2(new_n394), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n359), .B(new_n397), .C1(new_n400), .C2(new_n401), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT38), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n416), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n429), .A2(new_n432), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n483), .A2(KEYINPUT39), .A3(new_n433), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n439), .A2(new_n434), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT39), .B(new_n485), .C1(new_n483), .C2(new_n433), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n454), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT40), .A4(new_n454), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(new_n452), .A3(new_n417), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n389), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n389), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n459), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n267), .B1(new_n468), .B2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G183gat), .B(G211gat), .Z(new_n497));
  XNOR2_X1  g296(.A(G127gat), .B(G155gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G64gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT91), .ZN(new_n502));
  INV_X1    g301(.A(G57gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(G64gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(G64gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT9), .ZN(new_n508));
  NAND2_X1  g307(.A1(G71gat), .A2(G78gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n500), .A2(G57gat), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT9), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(new_n507), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n506), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT93), .ZN(new_n518));
  AND2_X1   g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n499), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n518), .A2(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n498), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n522), .B2(new_n525), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n208), .A2(new_n209), .B1(KEYINPUT21), .B2(new_n515), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n520), .A2(new_n521), .A3(new_n499), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n498), .B1(new_n523), .B2(new_n524), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n497), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n532), .A3(new_n536), .ZN(new_n540));
  INV_X1    g339(.A(new_n497), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G134gat), .B(G162gat), .Z(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT95), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G92gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT8), .ZN(new_n550));
  AND2_X1   g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n549), .A2(G85gat), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT94), .ZN(new_n553));
  OAI211_X1 g352(.A(G85gat), .B(G92gat), .C1(new_n553), .C2(KEYINPUT7), .ZN(new_n554));
  NAND2_X1  g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT7), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT94), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n554), .A2(new_n557), .B1(new_n553), .B2(KEYINPUT7), .ZN(new_n558));
  NOR2_X1   g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n552), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n557), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n550), .B1(G99gat), .B2(G106gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT95), .B(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n562), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n230), .B2(new_n233), .ZN(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n571), .A2(new_n236), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n580), .B2(new_n582), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n544), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  INV_X1    g388(.A(new_n544), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n506), .A2(new_n510), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n512), .A2(new_n514), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n561), .B2(new_n570), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n560), .B1(new_n552), .B2(new_n558), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n565), .A2(new_n562), .A3(new_n569), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n515), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n571), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n595), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n595), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT98), .ZN(new_n612));
  XOR2_X1   g411(.A(G176gat), .B(G204gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n607), .A2(new_n609), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n496), .A2(new_n543), .A3(new_n593), .A4(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n472), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(G1gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(G1324gat));
  INV_X1    g422(.A(new_n417), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(KEYINPUT100), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(G8gat), .ZN(new_n630));
  OAI221_X1 g429(.A(new_n627), .B1(KEYINPUT42), .B2(new_n626), .C1(new_n628), .C2(new_n630), .ZN(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n620), .B2(new_n471), .ZN(new_n632));
  INV_X1    g431(.A(new_n470), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(G15gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n620), .B2(new_n634), .ZN(G1326gat));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n389), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT43), .B(G22gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(new_n543), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n592), .A3(new_n619), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n496), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n642), .A2(G29gat), .A3(new_n472), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT45), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n494), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n459), .A2(new_n493), .A3(KEYINPUT103), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n471), .A2(new_n492), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n468), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n592), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n468), .A2(new_n495), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n593), .A2(new_n656), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n655), .A2(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n543), .A2(new_n267), .A3(new_n618), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G29gat), .B1(new_n661), .B2(new_n472), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n645), .A2(KEYINPUT45), .A3(new_n646), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n649), .A2(new_n662), .A3(new_n663), .ZN(G1328gat));
  OAI21_X1  g463(.A(G36gat), .B1(new_n661), .B2(new_n624), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n642), .A2(G36gat), .A3(new_n624), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n667), .A2(KEYINPUT46), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT46), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(G1329gat));
  NOR3_X1   g470(.A1(new_n642), .A2(G43gat), .A3(new_n633), .ZN(new_n672));
  INV_X1    g471(.A(new_n471), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n659), .A2(new_n673), .A3(new_n660), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n674), .B2(G43gat), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n675), .A2(KEYINPUT105), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n675), .B2(KEYINPUT105), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(G1330gat));
  NAND2_X1  g479(.A1(new_n493), .A2(G50gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n642), .A2(new_n389), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n661), .A2(new_n681), .B1(G50gat), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g483(.A1(new_n543), .A2(new_n267), .A3(new_n593), .A4(new_n618), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n468), .B2(new_n653), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n473), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g487(.A(new_n624), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n690), .B(new_n691), .Z(G1333gat));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n673), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n633), .A2(G71gat), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n693), .A2(G71gat), .B1(new_n686), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1334gat));
  NAND2_X1  g496(.A1(new_n686), .A2(new_n493), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g498(.A1(new_n393), .A2(new_n459), .A3(KEYINPUT35), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT86), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT35), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n471), .A2(new_n492), .A3(new_n494), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n658), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n543), .A2(new_n266), .A3(new_n619), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n593), .B1(new_n468), .B2(new_n653), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(KEYINPUT44), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n568), .A3(new_n472), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n543), .A2(new_n266), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n654), .A2(new_n592), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n619), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n473), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n710), .B1(new_n717), .B2(new_n568), .ZN(G1336gat));
  NOR2_X1   g517(.A1(new_n709), .A2(new_n624), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n709), .A2(KEYINPUT109), .A3(new_n624), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n549), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n714), .A2(new_n715), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n725), .A2(new_n545), .A3(new_n417), .A4(new_n618), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n719), .A2(new_n567), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT108), .B(new_n549), .C1(new_n709), .C2(new_n624), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT52), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(G1337gat));
  INV_X1    g532(.A(G99gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n709), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n673), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(KEYINPUT110), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT110), .B2(new_n736), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n716), .A2(new_n734), .A3(new_n470), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1338gat));
  NOR3_X1   g539(.A1(new_n389), .A2(G106gat), .A3(new_n619), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT111), .ZN(new_n742));
  AND4_X1   g541(.A1(KEYINPUT51), .A2(new_n654), .A3(new_n592), .A4(new_n711), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT51), .B1(new_n708), .B2(new_n711), .ZN(new_n744));
  OAI211_X1 g543(.A(KEYINPUT112), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G106gat), .B1(new_n709), .B2(new_n389), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT112), .B1(new_n725), .B2(new_n742), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT53), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT113), .B(KEYINPUT53), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n735), .B2(new_n493), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n709), .A2(KEYINPUT114), .A3(new_n389), .ZN(new_n755));
  OAI21_X1  g554(.A(G106gat), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT53), .B1(new_n725), .B2(new_n741), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n751), .A2(new_n752), .A3(new_n758), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n604), .A2(new_n605), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n594), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n614), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n604), .A2(new_n605), .A3(new_n595), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT115), .A4(new_n595), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n606), .A2(new_n762), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n617), .B1(new_n771), .B2(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  INV_X1    g572(.A(new_n764), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(KEYINPUT55), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n760), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n780), .A2(KEYINPUT116), .A3(new_n617), .A4(new_n775), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n266), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n261), .A2(new_n257), .ZN(new_n783));
  INV_X1    g582(.A(new_n245), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n243), .A2(new_n237), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n243), .A2(new_n787), .A3(new_n237), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n235), .B1(new_n234), .B2(new_n237), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n783), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n618), .A2(new_n265), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n592), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n265), .A2(new_n791), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n592), .A3(new_n781), .A4(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n639), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n543), .A2(new_n267), .A3(new_n593), .A4(new_n619), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT118), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n472), .A2(new_n417), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n393), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(G113gat), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n806), .A2(new_n807), .A3(new_n267), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n335), .A2(new_n463), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n803), .A2(new_n809), .A3(new_n493), .ZN(new_n810));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810), .B2(new_n266), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n808), .A2(new_n811), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n806), .B2(new_n619), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT119), .ZN(new_n814));
  INV_X1    g613(.A(G120gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n810), .A2(new_n815), .A3(new_n618), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n806), .B2(new_n639), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n810), .A2(new_n300), .A3(new_n543), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n809), .A2(new_n493), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n304), .A3(new_n821), .A4(new_n592), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT56), .Z(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n806), .B2(new_n593), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(G1343gat));
  NAND2_X1  g624(.A1(new_n471), .A2(new_n493), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n803), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n267), .A2(G141gat), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT58), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n493), .A2(KEYINPUT57), .ZN(new_n830));
  AND4_X1   g629(.A1(new_n267), .A2(new_n543), .A3(new_n593), .A4(new_n619), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n792), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n266), .A2(new_n617), .A3(new_n775), .A4(new_n780), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n592), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n639), .B1(new_n835), .B2(new_n796), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n831), .B1(KEYINPUT122), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n639), .C1(new_n835), .C2(new_n796), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n830), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n797), .A2(new_n798), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n798), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n493), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n471), .A2(new_n802), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n847), .A2(new_n267), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(G141gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n829), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n827), .A2(new_n828), .ZN(new_n852));
  INV_X1    g651(.A(new_n840), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n799), .A2(new_n800), .A3(new_n389), .ZN(new_n854));
  INV_X1    g653(.A(new_n846), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n848), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(KEYINPUT123), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n847), .B2(new_n848), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n860), .A3(new_n266), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n852), .B1(new_n861), .B2(G141gat), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n851), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n851), .B(KEYINPUT124), .C1(new_n862), .C2(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1344gat));
  INV_X1    g667(.A(G148gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n827), .A2(new_n869), .A3(new_n618), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n858), .A2(new_n860), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n619), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(KEYINPUT59), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n592), .A2(new_n794), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n776), .A3(new_n772), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n835), .A2(new_n875), .A3(KEYINPUT125), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n543), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n835), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n389), .B1(new_n879), .B2(new_n798), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .B1(new_n845), .B2(new_n846), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n618), .ZN(new_n882));
  OAI21_X1  g681(.A(G148gat), .B1(new_n882), .B2(new_n848), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n870), .B1(new_n873), .B2(new_n884), .ZN(G1345gat));
  OAI21_X1  g684(.A(G155gat), .B1(new_n871), .B2(new_n639), .ZN(new_n886));
  INV_X1    g685(.A(new_n827), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n639), .A2(G155gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n871), .B2(new_n593), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n593), .A2(G162gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n887), .B2(new_n891), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n473), .A2(new_n624), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n801), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(new_n821), .ZN(new_n895));
  AOI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n266), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n805), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n274), .A3(new_n267), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(G1348gat));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n275), .A3(new_n618), .ZN(new_n900));
  OAI21_X1  g699(.A(G176gat), .B1(new_n897), .B2(new_n619), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1349gat));
  NOR2_X1   g701(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n895), .A2(new_n284), .A3(new_n543), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n897), .B2(new_n639), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n906), .B(new_n907), .Z(G1350gat));
  NAND3_X1  g707(.A1(new_n895), .A2(new_n285), .A3(new_n592), .ZN(new_n909));
  OAI21_X1  g708(.A(G190gat), .B1(new_n897), .B2(new_n593), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT127), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n911), .B2(KEYINPUT127), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n909), .B1(new_n912), .B2(new_n914), .ZN(G1351gat));
  INV_X1    g714(.A(new_n826), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n266), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n881), .A2(new_n471), .A3(new_n893), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n266), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g721(.A1(new_n917), .A2(G204gat), .A3(new_n619), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n471), .A2(new_n893), .ZN(new_n925));
  OAI21_X1  g724(.A(G204gat), .B1(new_n882), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1353gat));
  AOI21_X1  g726(.A(new_n354), .B1(new_n920), .B2(new_n543), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT63), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n354), .A3(new_n543), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1354gat));
  NAND3_X1  g730(.A1(new_n918), .A2(new_n355), .A3(new_n592), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n920), .A2(new_n592), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n355), .ZN(G1355gat));
endmodule


