//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G15gat), .A2(G22gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G15gat), .A2(G22gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n211), .A2(new_n212), .A3(G1gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n214), .A3(G8gat), .ZN(new_n215));
  INV_X1    g014(.A(G8gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n208), .B(new_n213), .C1(new_n209), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  AND2_X1   g018(.A1(G71gat), .A2(G78gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G57gat), .B(G64gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G57gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G64gat), .ZN(new_n227));
  INV_X1    g026(.A(G64gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G57gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G71gat), .B(G78gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n224), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT93), .ZN(new_n236));
  INV_X1    g035(.A(G231gat), .ZN(new_n237));
  INV_X1    g036(.A(G233gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT93), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n235), .B(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n237), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n219), .ZN(new_n244));
  XOR2_X1   g043(.A(G127gat), .B(G155gat), .Z(new_n245));
  XOR2_X1   g044(.A(new_n244), .B(new_n245), .Z(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n239), .B2(new_n243), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n205), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n239), .A2(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n246), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n204), .A3(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(G232gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT41), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G43gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(G50gat), .ZN(new_n261));
  INV_X1    g060(.A(G50gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(G43gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT14), .ZN(new_n265));
  INV_X1    g064(.A(G29gat), .ZN(new_n266));
  INV_X1    g065(.A(G36gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n266), .A2(new_n267), .ZN(new_n271));
  OAI211_X1 g070(.A(KEYINPUT15), .B(new_n264), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT15), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n261), .B2(new_n263), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n262), .A2(G43gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n260), .A2(G50gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT15), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(new_n269), .ZN(new_n278));
  INV_X1    g077(.A(new_n271), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G99gat), .A2(G106gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g082(.A1(G85gat), .A2(G92gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT7), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G85gat), .ZN(new_n287));
  INV_X1    g086(.A(G92gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n283), .A2(new_n286), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G99gat), .B(G106gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g096(.A1(KEYINPUT8), .A2(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n259), .B1(new_n281), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n302), .B(new_n305), .C1(new_n272), .C2(new_n280), .ZN(new_n306));
  AND4_X1   g105(.A1(new_n303), .A2(new_n272), .A3(new_n304), .A4(new_n280), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n256), .B(new_n301), .C1(new_n308), .C2(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(new_n302), .ZN(new_n310));
  INV_X1    g109(.A(new_n305), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n281), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n272), .A2(new_n280), .A3(new_n303), .A4(new_n304), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n300), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n301), .ZN(new_n315));
  OAI21_X1  g114(.A(G190gat), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n316), .A3(G218gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(G218gat), .B1(new_n309), .B2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n257), .A2(new_n258), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n321), .B(KEYINPUT94), .Z(new_n322));
  XNOR2_X1  g121(.A(G134gat), .B(G162gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OR3_X1    g124(.A1(new_n319), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n319), .B2(new_n320), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n255), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G15gat), .B(G43gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G71gat), .B(G99gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT69), .B(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(G183gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT70), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g139(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n342));
  NAND2_X1  g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(KEYINPUT68), .A3(new_n344), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n338), .A2(new_n340), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT66), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT23), .ZN(new_n353));
  NAND2_X1  g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT25), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n336), .A2(new_n256), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n345), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n351), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT67), .A2(KEYINPUT25), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n355), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT26), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n354), .B1(new_n352), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n371), .A2(KEYINPUT73), .B1(new_n370), .B2(new_n352), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(KEYINPUT73), .B2(new_n371), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n335), .A2(KEYINPUT28), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT72), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n376), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n374), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n335), .B2(new_n375), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n373), .B(new_n343), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n369), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G113gat), .B(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT1), .ZN(new_n385));
  XNOR2_X1  g184(.A(G127gat), .B(G134gat), .ZN(new_n386));
  OR2_X1    g185(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n387), .B(new_n386), .C1(new_n384), .C2(KEYINPUT1), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT64), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n365), .B1(new_n348), .B2(new_n358), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(new_n368), .ZN(new_n396));
  INV_X1    g195(.A(new_n391), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n382), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n334), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n394), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n396), .A2(new_n397), .A3(new_n382), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n396), .B2(new_n382), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT75), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT34), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n401), .A2(new_n409), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(KEYINPUT34), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n399), .B2(KEYINPUT32), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n399), .A2(KEYINPUT32), .A3(new_n412), .ZN(new_n414));
  OAI22_X1  g213(.A1(new_n410), .A2(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n401), .A2(new_n409), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n414), .A2(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n409), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G78gat), .B(G106gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT31), .B(G50gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G22gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT84), .ZN(new_n426));
  NAND2_X1  g225(.A1(G228gat), .A2(G233gat), .ZN(new_n427));
  XOR2_X1   g226(.A(G155gat), .B(G162gat), .Z(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT77), .B(G162gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G155gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n430), .B2(KEYINPUT2), .ZN(new_n431));
  INV_X1    g230(.A(G141gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G148gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT76), .B(G148gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT2), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n432), .A2(G148gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n428), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT78), .B1(new_n442), .B2(KEYINPUT3), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n431), .A2(new_n435), .B1(new_n440), .B2(new_n428), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G197gat), .B(G204gat), .ZN(new_n449));
  INV_X1    g248(.A(G211gat), .ZN(new_n450));
  INV_X1    g249(.A(G218gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n449), .B1(KEYINPUT22), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G211gat), .B(G218gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n436), .A2(KEYINPUT79), .A3(new_n441), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT79), .B1(new_n436), .B2(new_n441), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n446), .B1(new_n455), .B2(KEYINPUT29), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n448), .A2(new_n456), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n427), .B1(new_n460), .B2(new_n442), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n448), .B2(new_n456), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n427), .A2(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT83), .B(new_n463), .C1(new_n448), .C2(new_n456), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n426), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n427), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  AND4_X1   g269(.A1(new_n426), .A2(new_n469), .A3(new_n470), .A4(new_n467), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n425), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n470), .A3(new_n467), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT84), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n466), .A2(new_n426), .A3(new_n467), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n424), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n420), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n391), .C1(new_n457), .C2(new_n458), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n436), .A2(new_n391), .A3(new_n441), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n444), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n479), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n391), .B1(new_n442), .B2(KEYINPUT3), .ZN(new_n489));
  INV_X1    g288(.A(new_n447), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT80), .B1(new_n444), .B2(new_n391), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(KEYINPUT82), .A3(new_n481), .ZN(new_n496));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n488), .A2(new_n492), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n480), .B1(new_n493), .B2(new_n494), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT4), .B(new_n391), .C1(new_n457), .C2(new_n458), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n492), .A2(new_n501), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT81), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n485), .A2(new_n486), .B1(new_n442), .B2(new_n397), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n497), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n493), .A2(new_n494), .B1(new_n444), .B2(new_n391), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT81), .A3(new_n498), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n503), .A2(new_n506), .A3(new_n508), .A4(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(new_n287), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT0), .B(G57gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516));
  INV_X1    g315(.A(new_n514), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI211_X1 g318(.A(new_n516), .B(new_n517), .C1(new_n500), .C2(new_n509), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G226gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n238), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT29), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n383), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n396), .B2(new_n382), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n455), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n383), .A2(new_n523), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n396), .B2(new_n382), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n456), .C1(new_n530), .C2(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G8gat), .B(G36gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(G64gat), .B(G92gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  OR3_X1    g334(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n535), .ZN(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n538), .A3(new_n531), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(KEYINPUT30), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n519), .A2(new_n521), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n478), .A2(KEYINPUT87), .A3(KEYINPUT35), .A4(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n415), .A2(new_n419), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n476), .A4(new_n472), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n519), .A2(new_n521), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n536), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n543), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n518), .A2(new_n516), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n517), .B1(new_n500), .B2(new_n509), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(new_n520), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n528), .A2(new_n555), .A3(new_n531), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n528), .A2(new_n555), .A3(new_n531), .A4(KEYINPUT37), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT38), .B1(new_n560), .B2(new_n538), .ZN(new_n561));
  INV_X1    g360(.A(new_n539), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n538), .B1(new_n558), .B2(new_n559), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT38), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n554), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n488), .A2(new_n492), .A3(new_n496), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT39), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n498), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n517), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT39), .B1(new_n507), .B2(new_n498), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n567), .B2(new_n498), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT85), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT40), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575));
  OAI211_X1 g374(.A(KEYINPUT85), .B(new_n575), .C1(new_n570), .C2(new_n572), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n540), .A2(new_n536), .A3(new_n515), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n477), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n566), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n544), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT36), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n548), .A2(new_n477), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n330), .B1(new_n550), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n218), .B1(new_n306), .B2(new_n307), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n215), .A2(new_n217), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n281), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n588), .A2(KEYINPUT18), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(KEYINPUT13), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n590), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n589), .A2(new_n281), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n592), .A2(new_n597), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT91), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n588), .A2(new_n612), .A3(new_n590), .A4(new_n591), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n606), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT18), .B1(new_n609), .B2(KEYINPUT91), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n607), .B1(new_n616), .B2(new_n613), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n606), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n234), .B1(new_n294), .B2(new_n299), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n291), .A2(new_n293), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n297), .A2(new_n292), .A3(new_n298), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n225), .A3(new_n623), .A4(new_n233), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n300), .A2(KEYINPUT10), .A3(new_n225), .A4(new_n233), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n620), .A2(new_n624), .ZN(new_n630));
  INV_X1    g429(.A(new_n628), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n633), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n587), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n546), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT96), .B(G1gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1324gat));
  INV_X1    g444(.A(new_n642), .ZN(new_n646));
  INV_X1    g445(.A(new_n547), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(G8gat), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(KEYINPUT42), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(KEYINPUT97), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n651), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n657), .A3(new_n584), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n646), .A2(new_n544), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(G1326gat));
  OR3_X1    g459(.A1(new_n642), .A2(KEYINPUT98), .A3(new_n579), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT98), .B1(new_n642), .B2(new_n579), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  AOI21_X1  g464(.A(new_n329), .B1(new_n550), .B2(new_n586), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n255), .A2(new_n619), .A3(new_n640), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n554), .A2(new_n266), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n668), .A2(KEYINPUT99), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT99), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(KEYINPUT45), .A3(new_n671), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n255), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n251), .A2(KEYINPUT100), .A3(new_n254), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n641), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n566), .A2(new_n578), .A3(new_n579), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n583), .B(new_n582), .C1(new_n579), .C2(new_n541), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n549), .B(new_n542), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n685), .B2(new_n328), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n682), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n681), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(KEYINPUT101), .A3(new_n554), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G29gat), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n689), .B2(new_n554), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n674), .B(new_n675), .C1(new_n691), .C2(new_n692), .ZN(G1328gat));
  NOR3_X1   g492(.A1(new_n668), .A2(G36gat), .A3(new_n547), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT46), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n689), .A2(new_n647), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n267), .B2(new_n696), .ZN(G1329gat));
  NOR2_X1   g496(.A1(new_n584), .A2(new_n260), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n260), .B1(new_n668), .B2(new_n420), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1330gat));
  AOI21_X1  g503(.A(new_n262), .B1(new_n689), .B2(new_n477), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n666), .A2(new_n262), .A3(new_n477), .A4(new_n667), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n705), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1331gat));
  XNOR2_X1  g510(.A(new_n617), .B(new_n606), .ZN(new_n712));
  INV_X1    g511(.A(new_n640), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n587), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n546), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(new_n226), .ZN(G1332gat));
  INV_X1    g516(.A(KEYINPUT49), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n647), .B1(new_n718), .B2(new_n228), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n715), .A2(KEYINPUT103), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT103), .B1(new_n715), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n228), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n715), .B2(new_n584), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n420), .A2(G71gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n715), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g527(.A1(new_n715), .A2(new_n579), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT104), .B(G78gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n255), .A2(new_n712), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n563), .A2(new_n564), .ZN(new_n733));
  AOI211_X1 g532(.A(KEYINPUT38), .B(new_n538), .C1(new_n558), .C2(new_n559), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n733), .A2(new_n734), .A3(new_n562), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n477), .B1(new_n735), .B2(new_n554), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n684), .B1(new_n736), .B2(new_n578), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n542), .A2(new_n549), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n328), .B(new_n732), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n713), .B1(new_n739), .B2(KEYINPUT51), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n685), .A2(new_n741), .A3(new_n328), .A4(new_n732), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n287), .A3(new_n554), .ZN(new_n744));
  INV_X1    g543(.A(new_n255), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n714), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  AOI211_X1 g546(.A(KEYINPUT44), .B(new_n329), .C1(new_n550), .C2(new_n586), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n686), .ZN(new_n749));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749), .B2(new_n546), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n750), .ZN(G1336gat));
  OAI211_X1 g550(.A(new_n647), .B(new_n747), .C1(new_n748), .C2(new_n686), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(new_n753), .A3(G92gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT51), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n547), .A2(G92gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n640), .A3(new_n742), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(new_n757), .C1(new_n758), .C2(new_n753), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n752), .A2(new_n760), .A3(G92gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n752), .B2(G92gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n757), .A2(new_n758), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n759), .B1(new_n764), .B2(new_n753), .ZN(G1337gat));
  XOR2_X1   g564(.A(KEYINPUT108), .B(G99gat), .Z(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n743), .A2(new_n544), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n749), .B2(new_n584), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1338gat));
  NOR2_X1   g569(.A1(new_n579), .A2(G106gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n740), .A2(new_n742), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n477), .B(new_n747), .C1(new_n748), .C2(new_n686), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n740), .A2(KEYINPUT109), .A3(new_n742), .A4(new_n771), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT53), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n775), .B2(G106gat), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT110), .A3(new_n772), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT110), .B1(new_n780), .B2(new_n772), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(new_n605), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n614), .A2(new_n608), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n591), .B1(new_n588), .B2(new_n590), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n595), .A2(new_n596), .A3(new_n594), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n604), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n640), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n790));
  AND4_X1   g589(.A1(KEYINPUT111), .A2(new_n629), .A3(KEYINPUT54), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n627), .B2(new_n628), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT111), .B1(new_n793), .B2(new_n790), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n795));
  INV_X1    g594(.A(new_n636), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n631), .B1(new_n625), .B2(new_n626), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n792), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n627), .A2(new_n792), .A3(new_n628), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT112), .B1(new_n799), .B2(new_n636), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n791), .A2(new_n794), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT54), .B(new_n631), .C1(new_n625), .C2(new_n626), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n795), .B1(new_n804), .B2(new_n796), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n636), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(KEYINPUT55), .C1(new_n794), .C2(new_n791), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n638), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n789), .B1(new_n619), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n637), .B1(new_n801), .B2(new_n802), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n808), .C1(new_n615), .C2(new_n618), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n789), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n811), .A2(new_n329), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n629), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n793), .A2(KEYINPUT111), .A3(new_n790), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n819), .A2(new_n820), .B1(new_n805), .B2(new_n806), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n638), .B1(new_n821), .B2(KEYINPUT55), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n801), .A2(new_n802), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n785), .A2(new_n788), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n328), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n824), .A2(new_n328), .A3(new_n828), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n679), .B1(new_n816), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n255), .A2(new_n619), .A3(new_n713), .A4(new_n329), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n478), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n546), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n547), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT115), .ZN(new_n840));
  INV_X1    g639(.A(G113gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n712), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n839), .B2(new_n619), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1340gat));
  INV_X1    g643(.A(G120gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(new_n845), .A3(new_n640), .ZN(new_n846));
  OAI21_X1  g645(.A(G120gat), .B1(new_n839), .B2(new_n713), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n839), .A2(new_n851), .A3(new_n680), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n255), .A3(new_n547), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(G1342gat));
  NAND2_X1  g653(.A1(new_n547), .A2(new_n328), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT117), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n837), .A2(G134gat), .A3(new_n856), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT56), .Z(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n839), .B2(new_n329), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n477), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n584), .A2(new_n554), .A3(new_n547), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n712), .A2(new_n432), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(KEYINPUT58), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n871));
  AOI21_X1  g670(.A(new_n871), .B1(new_n834), .B2(new_n477), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873));
  INV_X1    g672(.A(new_n789), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n874), .B1(new_n824), .B2(new_n712), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n329), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n813), .A2(new_n876), .A3(new_n789), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n830), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n745), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n873), .B(new_n579), .C1(new_n880), .C2(new_n832), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n712), .B(new_n864), .C1(new_n872), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G141gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n870), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n882), .A2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n887), .B2(new_n869), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n881), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n863), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n640), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n477), .B(new_n871), .C1(new_n831), .C2(new_n833), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n826), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n328), .B1(new_n810), .B2(KEYINPUT119), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n875), .A2(new_n876), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n832), .B1(new_n899), .B2(new_n255), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n900), .B2(new_n477), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n713), .A3(new_n863), .ZN(new_n903));
  NAND2_X1  g702(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n865), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n892), .B1(new_n905), .B2(new_n640), .ZN(new_n906));
  OAI221_X1 g705(.A(new_n893), .B1(new_n903), .B2(new_n904), .C1(new_n906), .C2(new_n434), .ZN(G1345gat));
  AOI21_X1  g706(.A(G155gat), .B1(new_n905), .B2(new_n255), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n679), .A2(G155gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n891), .B2(new_n909), .ZN(G1346gat));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n328), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n429), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n856), .A2(new_n429), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n554), .A3(new_n584), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n861), .B2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n554), .A2(new_n547), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n916), .A2(new_n478), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n834), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n712), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n640), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g721(.A(new_n336), .B1(new_n918), .B2(new_n679), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n377), .A2(new_n378), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n255), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  NAND2_X1  g727(.A1(new_n918), .A2(new_n328), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G190gat), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(KEYINPUT123), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n934));
  INV_X1    g733(.A(new_n335), .ZN(new_n935));
  OAI22_X1  g734(.A1(new_n933), .A2(new_n934), .B1(new_n935), .B2(new_n929), .ZN(G1351gat));
  OR2_X1    g735(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n584), .A2(new_n916), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n619), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n862), .A2(new_n939), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n619), .A2(G197gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  OAI21_X1  g743(.A(G204gat), .B1(new_n940), .B2(new_n713), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n713), .A2(G204gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n862), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n947), .B2(KEYINPUT62), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n945), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(G1353gat));
  INV_X1    g751(.A(new_n942), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n450), .A3(new_n255), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n255), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n895), .B2(new_n901), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n957), .A2(KEYINPUT126), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n826), .B1(new_n877), .B2(new_n878), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n833), .B1(new_n960), .B2(new_n745), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n873), .B1(new_n961), .B2(new_n579), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n955), .B1(new_n962), .B2(new_n894), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n963), .B2(new_n450), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n876), .B1(new_n813), .B2(new_n789), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n878), .A2(new_n966), .A3(new_n328), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n745), .B1(new_n967), .B2(new_n896), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n579), .B1(new_n968), .B2(new_n832), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n894), .B1(new_n969), .B2(KEYINPUT57), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n450), .B1(new_n970), .B2(new_n956), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT126), .B1(new_n971), .B2(KEYINPUT63), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n954), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(KEYINPUT127), .B(new_n954), .C1(new_n965), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1354gat));
  NOR3_X1   g776(.A1(new_n940), .A2(new_n451), .A3(new_n329), .ZN(new_n978));
  AOI21_X1  g777(.A(G218gat), .B1(new_n953), .B2(new_n328), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


