

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U554 ( .A(KEYINPUT64), .B(n523), .ZN(n648) );
  INV_X4 U555 ( .A(G2105), .ZN(n604) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n685) );
  XNOR2_X2 U557 ( .A(n685), .B(KEYINPUT89), .ZN(n785) );
  AND2_X1 U558 ( .A1(n560), .A2(n559), .ZN(n562) );
  BUF_X1 U559 ( .A(n608), .Z(n519) );
  XNOR2_X1 U560 ( .A(n556), .B(n555), .ZN(n608) );
  XNOR2_X2 U561 ( .A(n562), .B(n561), .ZN(G160) );
  XOR2_X1 U562 ( .A(KEYINPUT76), .B(n569), .Z(n520) );
  AND2_X1 U563 ( .A1(n907), .A2(n698), .ZN(n699) );
  INV_X1 U564 ( .A(KEYINPUT96), .ZN(n690) );
  XNOR2_X1 U565 ( .A(KEYINPUT95), .B(KEYINPUT29), .ZN(n724) );
  XNOR2_X1 U566 ( .A(n725), .B(n724), .ZN(n728) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  AND2_X1 U568 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U569 ( .A(G120), .ZN(G236) );
  INV_X1 U570 ( .A(G69), .ZN(G235) );
  INV_X1 U571 ( .A(G132), .ZN(G219) );
  INV_X1 U572 ( .A(G82), .ZN(G220) );
  NOR2_X1 U573 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U574 ( .A1(G88), .A2(n639), .ZN(n522) );
  INV_X1 U575 ( .A(G651), .ZN(n525) );
  NOR2_X2 U576 ( .A1(n626), .A2(n525), .ZN(n644) );
  NAND2_X1 U577 ( .A1(G75), .A2(n644), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n626), .A2(G651), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n648), .A2(G50), .ZN(n524) );
  XNOR2_X1 U581 ( .A(n524), .B(KEYINPUT84), .ZN(n528) );
  NOR2_X1 U582 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X2 U583 ( .A(KEYINPUT1), .B(n526), .Z(n640) );
  NAND2_X1 U584 ( .A1(n640), .A2(G62), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(G166) );
  NAND2_X1 U587 ( .A1(G64), .A2(n640), .ZN(n532) );
  NAND2_X1 U588 ( .A1(G52), .A2(n648), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n537) );
  NAND2_X1 U590 ( .A1(G90), .A2(n639), .ZN(n534) );
  NAND2_X1 U591 ( .A1(G77), .A2(n644), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U593 ( .A(KEYINPUT9), .B(n535), .Z(n536) );
  NOR2_X1 U594 ( .A1(n537), .A2(n536), .ZN(G171) );
  NAND2_X1 U595 ( .A1(n639), .A2(G89), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT4), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G76), .A2(n644), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U599 ( .A(KEYINPUT5), .B(n541), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G63), .A2(n640), .ZN(n543) );
  NAND2_X1 U601 ( .A1(G51), .A2(n648), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n544) );
  XNOR2_X1 U604 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U606 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  XNOR2_X2 U607 ( .A(G2104), .B(KEYINPUT66), .ZN(n603) );
  AND2_X1 U608 ( .A1(n604), .A2(G101), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n603), .A2(n549), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT67), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT23), .ZN(n560) );
  NOR2_X4 U612 ( .A1(n604), .A2(n603), .ZN(n880) );
  NAND2_X1 U613 ( .A1(G125), .A2(n880), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G2104), .A2(G2105), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT68), .B(n552), .Z(n677) );
  NAND2_X1 U616 ( .A1(G113), .A2(n677), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n558) );
  XNOR2_X1 U618 ( .A(KEYINPUT69), .B(KEYINPUT17), .ZN(n556) );
  NOR2_X1 U619 ( .A1(G2105), .A2(G2104), .ZN(n555) );
  AND2_X1 U620 ( .A1(G137), .A2(n608), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U622 ( .A(KEYINPUT65), .ZN(n561) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n563), .B(KEYINPUT74), .ZN(n564) );
  XNOR2_X1 U626 ( .A(KEYINPUT10), .B(n564), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n831) );
  NAND2_X1 U628 ( .A1(n831), .A2(G567), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT11), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT75), .B(n566), .ZN(G234) );
  NAND2_X1 U631 ( .A1(G56), .A2(n640), .ZN(n567) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n567), .Z(n573) );
  NAND2_X1 U633 ( .A1(n639), .A2(G81), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT12), .B(n568), .Z(n570) );
  NAND2_X1 U635 ( .A1(n644), .A2(G68), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n520), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G43), .A2(n648), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n969) );
  INV_X1 U641 ( .A(G860), .ZN(n596) );
  OR2_X1 U642 ( .A1(n969), .A2(n596), .ZN(G153) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G79), .A2(n644), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G54), .A2(n648), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G66), .A2(n640), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G92), .A2(n639), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U651 ( .A(KEYINPUT77), .B(n580), .Z(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X2 U653 ( .A(KEYINPUT15), .B(n583), .Z(n907) );
  INV_X1 U654 ( .A(n907), .ZN(n952) );
  INV_X1 U655 ( .A(G868), .ZN(n659) );
  NAND2_X1 U656 ( .A1(n952), .A2(n659), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n640), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G53), .A2(n648), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G91), .A2(n639), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G78), .A2(n644), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U664 ( .A(KEYINPUT71), .B(n590), .Z(n591) );
  NOR2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT72), .B(n593), .Z(G299) );
  NOR2_X1 U667 ( .A1(G286), .A2(n659), .ZN(n595) );
  NOR2_X1 U668 ( .A1(G299), .A2(G868), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n597), .A2(n907), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G559), .A2(n659), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n907), .A2(n599), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT79), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n969), .A2(G868), .ZN(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(G282) );
  AND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n877) );
  NAND2_X1 U679 ( .A1(n877), .A2(G99), .ZN(n606) );
  BUF_X1 U680 ( .A(n677), .Z(n881) );
  NAND2_X1 U681 ( .A1(G111), .A2(n881), .ZN(n605) );
  NAND2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n880), .A2(G123), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G135), .A2(n519), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n987) );
  XNOR2_X1 U688 ( .A(n987), .B(G2096), .ZN(n614) );
  INV_X1 U689 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G67), .A2(n640), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G93), .A2(n639), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G80), .A2(n644), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G55), .A2(n648), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n660) );
  XNOR2_X1 U699 ( .A(n969), .B(KEYINPUT80), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n907), .A2(G559), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n623), .B(n622), .ZN(n656) );
  NOR2_X1 U702 ( .A1(n656), .A2(G860), .ZN(n624) );
  XOR2_X1 U703 ( .A(n660), .B(n624), .Z(G145) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT82), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n626), .A2(G87), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G49), .A2(n648), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U709 ( .A1(n640), .A2(n629), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G85), .A2(n639), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G72), .A2(n644), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U714 ( .A(KEYINPUT70), .B(n634), .Z(n638) );
  NAND2_X1 U715 ( .A1(n648), .A2(G47), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G60), .A2(n640), .ZN(n635) );
  AND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U719 ( .A1(n639), .A2(G86), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n640), .A2(G61), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U722 ( .A(KEYINPUT83), .B(n643), .Z(n647) );
  NAND2_X1 U723 ( .A1(G73), .A2(n644), .ZN(n645) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n645), .Z(n646) );
  NOR2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G48), .A2(n648), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(G288), .ZN(n655) );
  XNOR2_X1 U729 ( .A(G290), .B(n660), .ZN(n653) );
  XNOR2_X1 U730 ( .A(G166), .B(G299), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(G305), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n904) );
  XNOR2_X1 U734 ( .A(n904), .B(n656), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n657), .A2(G868), .ZN(n658) );
  XOR2_X1 U736 ( .A(KEYINPUT85), .B(n658), .Z(n662) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U745 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n667) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U748 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(G96), .A2(n669), .ZN(n837) );
  NAND2_X1 U750 ( .A1(n837), .A2(G2106), .ZN(n675) );
  NOR2_X1 U751 ( .A1(G235), .A2(G236), .ZN(n670) );
  XNOR2_X1 U752 ( .A(KEYINPUT86), .B(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n671), .A2(G108), .ZN(n672) );
  NOR2_X1 U754 ( .A1(n672), .A2(G237), .ZN(n673) );
  XNOR2_X1 U755 ( .A(n673), .B(KEYINPUT87), .ZN(n838) );
  NAND2_X1 U756 ( .A1(n838), .A2(G567), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n839) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U759 ( .A1(n839), .A2(n676), .ZN(n836) );
  NAND2_X1 U760 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U761 ( .A1(G114), .A2(n677), .ZN(n678) );
  XNOR2_X1 U762 ( .A(n678), .B(KEYINPUT88), .ZN(n680) );
  NAND2_X1 U763 ( .A1(G138), .A2(n519), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n684) );
  NAND2_X1 U765 ( .A1(G126), .A2(n880), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G102), .A2(n877), .ZN(n681) );
  NAND2_X1 U767 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U768 ( .A1(n684), .A2(n683), .ZN(G164) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n787) );
  AND2_X2 U771 ( .A1(n787), .A2(n785), .ZN(n735) );
  INV_X1 U772 ( .A(G8), .ZN(n740) );
  OR2_X1 U773 ( .A1(G1966), .A2(n740), .ZN(n686) );
  NOR2_X1 U774 ( .A1(n735), .A2(n686), .ZN(n732) );
  INV_X1 U775 ( .A(n735), .ZN(n697) );
  NOR2_X1 U776 ( .A1(n697), .A2(G2084), .ZN(n730) );
  NOR2_X1 U777 ( .A1(n732), .A2(n730), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G8), .A2(n687), .ZN(n688) );
  XNOR2_X1 U779 ( .A(n688), .B(KEYINPUT30), .ZN(n689) );
  NOR2_X1 U780 ( .A1(G168), .A2(n689), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n691), .B(n690), .ZN(n695) );
  XOR2_X1 U782 ( .A(KEYINPUT25), .B(G2078), .Z(n932) );
  INV_X1 U783 ( .A(n735), .ZN(n702) );
  NOR2_X1 U784 ( .A1(n932), .A2(n702), .ZN(n693) );
  NOR2_X1 U785 ( .A1(n735), .A2(G1961), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n726) );
  NAND2_X1 U787 ( .A1(n726), .A2(G301), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT31), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n697), .A2(G1341), .ZN(n708) );
  INV_X1 U791 ( .A(n969), .ZN(n698) );
  AND2_X1 U792 ( .A1(n708), .A2(n699), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n735), .A2(G1996), .ZN(n700) );
  XNOR2_X1 U794 ( .A(n700), .B(KEYINPUT26), .ZN(n710) );
  NAND2_X1 U795 ( .A1(n701), .A2(n710), .ZN(n706) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n702), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n735), .A2(G1348), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT94), .ZN(n713) );
  AND2_X1 U801 ( .A1(n708), .A2(n698), .ZN(n709) );
  AND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  OR2_X1 U803 ( .A1(n711), .A2(n907), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n718) );
  NAND2_X1 U805 ( .A1(n735), .A2(G2072), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  INV_X1 U807 ( .A(G1956), .ZN(n1016) );
  NOR2_X1 U808 ( .A1(n1016), .A2(n735), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n720) );
  INV_X1 U810 ( .A(G299), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U814 ( .A(n721), .B(KEYINPUT28), .Z(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n725) );
  OR2_X1 U816 ( .A1(G301), .A2(n726), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n743) );
  AND2_X1 U818 ( .A1(n741), .A2(n743), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT97), .ZN(n734) );
  AND2_X1 U820 ( .A1(G8), .A2(n730), .ZN(n731) );
  NOR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n734), .A2(n733), .ZN(n751) );
  OR2_X1 U823 ( .A1(n735), .A2(n740), .ZN(n769) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n769), .ZN(n737) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n702), .ZN(n736) );
  NOR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n744) );
  AND2_X1 U829 ( .A1(n741), .A2(n744), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n748) );
  INV_X1 U831 ( .A(n744), .ZN(n746) );
  AND2_X1 U832 ( .A1(G286), .A2(G8), .ZN(n745) );
  OR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U835 ( .A(n749), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n764) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n948) );
  NOR2_X1 U839 ( .A1(n752), .A2(n948), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n764), .A2(n753), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NAND2_X1 U842 ( .A1(n754), .A2(n950), .ZN(n755) );
  XNOR2_X1 U843 ( .A(n755), .B(KEYINPUT98), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n756), .A2(n769), .ZN(n757) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n757), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n948), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U847 ( .A1(n758), .A2(n769), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n957) );
  AND2_X1 U850 ( .A1(n761), .A2(n957), .ZN(n774) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n769), .A2(n765), .ZN(n772) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U856 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  XNOR2_X1 U857 ( .A(KEYINPUT92), .B(n767), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U859 ( .A(KEYINPUT93), .B(n770), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n790) );
  NAND2_X1 U862 ( .A1(n877), .A2(G104), .ZN(n775) );
  XNOR2_X1 U863 ( .A(n775), .B(KEYINPUT90), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G140), .A2(n519), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT34), .B(n778), .ZN(n783) );
  NAND2_X1 U867 ( .A1(n880), .A2(G128), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G116), .A2(n881), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U870 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U872 ( .A(KEYINPUT36), .B(n784), .Z(n889) );
  XOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .Z(n812) );
  AND2_X1 U874 ( .A1(n889), .A2(n812), .ZN(n994) );
  INV_X1 U875 ( .A(n785), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n826) );
  NAND2_X1 U877 ( .A1(n994), .A2(n826), .ZN(n813) );
  XNOR2_X1 U878 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U879 ( .A1(n826), .A2(n966), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n813), .A2(n788), .ZN(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n809) );
  NAND2_X1 U882 ( .A1(G105), .A2(n877), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n791), .B(KEYINPUT38), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G129), .A2(n880), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G141), .A2(n519), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G117), .A2(n881), .ZN(n794) );
  XNOR2_X1 U888 ( .A(KEYINPUT91), .B(n794), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n894) );
  NAND2_X1 U891 ( .A1(G1996), .A2(n894), .ZN(n806) );
  NAND2_X1 U892 ( .A1(n877), .A2(G95), .ZN(n800) );
  NAND2_X1 U893 ( .A1(G107), .A2(n881), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G119), .A2(n880), .ZN(n802) );
  NAND2_X1 U896 ( .A1(G131), .A2(n519), .ZN(n801) );
  NAND2_X1 U897 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n897) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n897), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n990) );
  NAND2_X1 U901 ( .A1(n826), .A2(n990), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n809), .A2(n814), .ZN(n808) );
  INV_X1 U903 ( .A(KEYINPUT99), .ZN(n807) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n809), .A2(KEYINPUT99), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n829) );
  NAND2_X1 U907 ( .A1(n990), .A2(KEYINPUT99), .ZN(n825) );
  NOR2_X1 U908 ( .A1(n889), .A2(n812), .ZN(n999) );
  INV_X1 U909 ( .A(n813), .ZN(n822) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n894), .ZN(n983) );
  INV_X1 U911 ( .A(n814), .ZN(n818) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n897), .ZN(n988) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n815) );
  XNOR2_X1 U914 ( .A(KEYINPUT100), .B(n815), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n988), .A2(n816), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n983), .A2(n819), .ZN(n820) );
  XOR2_X1 U918 ( .A(KEYINPUT39), .B(n820), .Z(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n999), .A2(n823), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n831), .ZN(G217) );
  INV_X1 U926 ( .A(G661), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G2), .A2(G15), .ZN(n832) );
  NOR2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U929 ( .A(KEYINPUT104), .B(n834), .Z(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U932 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n839), .ZN(G319) );
  XNOR2_X1 U938 ( .A(G1996), .B(KEYINPUT41), .ZN(n849) );
  XOR2_X1 U939 ( .A(G1991), .B(G1986), .Z(n841) );
  XNOR2_X1 U940 ( .A(G1981), .B(G1966), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U942 ( .A(G1961), .B(G1956), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1976), .B(G1971), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U945 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2474), .B(KEYINPUT108), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U949 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT106), .B(G2678), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2096), .B(G2100), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U958 ( .A(G2084), .B(G2078), .Z(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U960 ( .A1(n877), .A2(G100), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G112), .A2(n881), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U963 ( .A1(G124), .A2(n880), .ZN(n862) );
  XOR2_X1 U964 ( .A(KEYINPUT109), .B(n862), .Z(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G136), .A2(n519), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U969 ( .A1(n880), .A2(G130), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G118), .A2(n881), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n877), .A2(G106), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT110), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G142), .A2(n519), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(n873), .ZN(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT45), .B(n874), .ZN(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n893) );
  NAND2_X1 U979 ( .A1(G139), .A2(n519), .ZN(n879) );
  NAND2_X1 U980 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n880), .A2(G127), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G115), .A2(n881), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT112), .B(n884), .Z(n885) );
  XNOR2_X1 U986 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  NOR2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT113), .B(n888), .Z(n978) );
  XOR2_X1 U989 ( .A(G162), .B(n978), .Z(n891) );
  XNOR2_X1 U990 ( .A(G164), .B(n889), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n894), .B(n987), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n902) );
  XNOR2_X1 U995 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n897), .B(KEYINPUT46), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(G160), .B(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U1001 ( .A(G286), .B(n904), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n969), .B(n905), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n906), .B(KEYINPUT115), .Z(n909) );
  XNOR2_X1 U1004 ( .A(n907), .B(G171), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1007 ( .A(KEYINPUT103), .B(G2446), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2454), .B(G2451), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n913), .B(G2430), .Z(n915) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n919) );
  XOR2_X1 U1013 ( .A(KEYINPUT102), .B(G2435), .Z(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT101), .B(G2438), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1016 ( .A(n919), .B(n918), .Z(n921) );
  XNOR2_X1 U1017 ( .A(G2443), .B(G2427), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n921), .B(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n922), .A2(G14), .ZN(n928) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n928), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(G229), .A2(G227), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(n928), .ZN(G401) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n1033) );
  XOR2_X1 U1029 ( .A(G1991), .B(G25), .Z(n929) );
  NAND2_X1 U1030 ( .A1(n929), .A2(G28), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(G1996), .B(G32), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(G27), .B(n932), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1039 ( .A(n939), .B(KEYINPUT53), .Z(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT118), .ZN(n946) );
  XOR2_X1 U1044 ( .A(G2084), .B(KEYINPUT54), .Z(n944) );
  XNOR2_X1 U1045 ( .A(G34), .B(n944), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n1032) );
  OR2_X1 U1047 ( .A1(n1033), .A2(n1032), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(G11), .A2(n947), .ZN(n1006) );
  INV_X1 U1049 ( .A(n948), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(n951), .B(KEYINPUT123), .ZN(n956) );
  XOR2_X1 U1052 ( .A(G1971), .B(G166), .Z(n954) );
  XNOR2_X1 U1053 ( .A(n952), .B(G1348), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(n959), .B(KEYINPUT57), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n960) );
  XNOR2_X1 U1060 ( .A(n961), .B(n960), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(n1016), .B(G299), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(n964), .B(KEYINPUT122), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G301), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n969), .ZN(n970) );
  NOR2_X1 U1068 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT124), .ZN(n977) );
  XOR2_X1 U1071 ( .A(G16), .B(KEYINPUT119), .Z(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT56), .B(n975), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n1004) );
  XOR2_X1 U1074 ( .A(G2072), .B(n978), .Z(n980) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1077 ( .A(KEYINPUT50), .B(n981), .Z(n986) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(KEYINPUT51), .B(n984), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n997) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G160), .B(G2084), .Z(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT116), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1033), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1038) );
  XNOR2_X1 U1095 ( .A(G1986), .B(G24), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT126), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G1966), .B(G21), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1027) );
  XOR2_X1 U1105 ( .A(G1981), .B(G6), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(n1016), .B(G20), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(G1341), .B(G19), .Z(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n1019) );
  XNOR2_X1 U1110 ( .A(G4), .B(n1019), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(n1020), .B(G1348), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1114 ( .A(n1025), .B(KEYINPUT60), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G5), .B(G1961), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1030), .Z(n1031) );
  NOR2_X1 U1119 ( .A1(G16), .A2(n1031), .ZN(n1036) );
  NAND2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(G29), .A2(n1034), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

