//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT79), .Z(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n193), .A2(KEYINPUT1), .A3(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n192), .A3(new_n194), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n204), .A3(new_n205), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT81), .B(G224), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n200), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n200), .B2(new_n208), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n217), .B2(KEYINPUT7), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G104), .B(G107), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT77), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(G107), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n221), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(G104), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n223), .A2(G107), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(G101), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n222), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n237));
  INV_X1    g051(.A(G113), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT2), .A2(G113), .ZN(new_n242));
  AND4_X1   g056(.A1(new_n236), .A2(new_n239), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT80), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n236), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n238), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G116), .B(G119), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n243), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT82), .B1(new_n234), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n243), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n234), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n239), .A3(new_n242), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n236), .A2(new_n241), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n248), .ZN(new_n261));
  OAI21_X1  g075(.A(G113), .B1(new_n252), .B2(new_n236), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT82), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n222), .A2(new_n229), .A3(new_n233), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G122), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT8), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n267), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT83), .B1(new_n267), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n219), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n234), .A2(new_n254), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G101), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n239), .A2(new_n242), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n260), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT4), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n281), .A3(G101), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n277), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n272), .A2(new_n273), .B1(new_n268), .B2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n219), .B(KEYINPUT84), .C1(new_n270), .C2(new_n271), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n190), .B(G902), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n272), .A2(new_n273), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(new_n268), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT85), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n289), .A2(KEYINPUT6), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n284), .A2(new_n268), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g110(.A(new_n217), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n189), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n267), .A2(new_n269), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n267), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n218), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n289), .B1(new_n304), .B2(KEYINPUT84), .ZN(new_n305));
  INV_X1    g119(.A(new_n286), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n291), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n190), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n290), .A2(KEYINPUT85), .A3(new_n291), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n189), .A3(new_n298), .A4(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n188), .B1(new_n299), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT86), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(KEYINPUT86), .B(new_n188), .C1(new_n299), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G234), .ZN(new_n317));
  OAI21_X1  g131(.A(G217), .B1(new_n317), .B2(G902), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT72), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n235), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n202), .A2(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n323), .A2(KEYINPUT73), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(KEYINPUT73), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT24), .B(G110), .Z(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G110), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n336), .A2(KEYINPUT16), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(G146), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(G146), .B1(new_n334), .B2(new_n337), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n327), .B(new_n332), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n191), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n338), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n346), .A2(KEYINPUT74), .A3(new_n332), .A4(new_n327), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n324), .A2(new_n325), .ZN(new_n349));
  OAI22_X1  g163(.A1(new_n349), .A2(new_n326), .B1(G110), .B2(new_n331), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n204), .A2(G140), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n336), .A2(new_n351), .A3(KEYINPUT75), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT75), .B1(new_n336), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n191), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n338), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT22), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(G137), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n348), .A2(new_n355), .A3(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n291), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(KEYINPUT25), .A3(new_n291), .A4(new_n362), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n320), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n361), .A2(new_n362), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n319), .A2(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT31), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT11), .ZN(new_n373));
  INV_X1    g187(.A(G134), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(G137), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(G137), .ZN(new_n376));
  INV_X1    g190(.A(G137), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(KEYINPUT11), .A3(G134), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G131), .ZN(new_n380));
  INV_X1    g194(.A(G131), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n375), .A2(new_n378), .A3(new_n381), .A4(new_n376), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n199), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n280), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n207), .B(new_n205), .C1(G128), .C2(new_n197), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n374), .B2(G137), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n377), .A2(KEYINPUT64), .A3(G134), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n376), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n382), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n386), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(KEYINPUT65), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(KEYINPUT65), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n387), .A2(new_n382), .A3(new_n392), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n199), .B1(new_n380), .B2(new_n382), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n385), .A2(KEYINPUT65), .A3(new_n393), .A4(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n395), .B1(new_n403), .B2(new_n280), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT26), .B(G101), .ZN(new_n405));
  NOR2_X1   g219(.A1(G237), .A2(G953), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G210), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n372), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n386), .B1(new_n401), .B2(new_n402), .ZN(new_n413));
  NOR4_X1   g227(.A1(new_n413), .A2(KEYINPUT31), .A3(new_n395), .A4(new_n410), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n395), .A2(KEYINPUT28), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n385), .A2(new_n393), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n280), .ZN(new_n420));
  AOI211_X1 g234(.A(KEYINPUT67), .B(new_n386), .C1(new_n385), .C2(new_n393), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n394), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n417), .B1(new_n422), .B2(KEYINPUT28), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n416), .B1(new_n423), .B2(new_n411), .ZN(new_n424));
  INV_X1    g238(.A(new_n417), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n280), .B1(new_n399), .B2(new_n400), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT67), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n386), .B1(new_n385), .B2(new_n393), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n418), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n395), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT28), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT68), .A3(new_n410), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(G472), .A2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT69), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT32), .B1(new_n434), .B2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n434), .A2(KEYINPUT32), .A3(new_n435), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n434), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n435), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n439), .A2(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT70), .B1(new_n432), .B2(new_n410), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n449));
  INV_X1    g263(.A(new_n404), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n410), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n423), .A2(new_n452), .A3(new_n411), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n449), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n395), .A2(new_n428), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n417), .B1(new_n456), .B2(KEYINPUT28), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n410), .A2(new_n449), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G472), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n371), .B1(new_n447), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  INV_X1    g277(.A(G227), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(KEYINPUT76), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(G110), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(G140), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n387), .A2(new_n229), .A3(new_n233), .A4(new_n222), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT10), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n387), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n277), .A2(new_n384), .A3(new_n282), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n383), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n206), .A2(new_n192), .A3(new_n194), .ZN(new_n476));
  AOI21_X1  g290(.A(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n477));
  INV_X1    g291(.A(new_n205), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n265), .A2(new_n479), .A3(KEYINPUT78), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n469), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT78), .B1(new_n265), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n383), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT12), .B(new_n383), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n468), .B(new_n475), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n468), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n474), .A2(new_n383), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n474), .A2(new_n383), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n463), .B(new_n291), .C1(new_n487), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G469), .A2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n488), .A3(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n475), .B1(new_n485), .B2(new_n486), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(new_n488), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n492), .B(new_n493), .C1(new_n463), .C2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT9), .B(G234), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G221), .B1(new_n499), .B2(G902), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(G113), .B(G122), .Z(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT93), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n223), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G237), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n213), .A3(G214), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT87), .A3(G143), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n193), .ZN(new_n510));
  NAND2_X1  g324(.A1(KEYINPUT87), .A2(G143), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n510), .A2(G214), .A3(new_n406), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n381), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(KEYINPUT17), .ZN(new_n515));
  INV_X1    g329(.A(new_n346), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n381), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n333), .A2(new_n191), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n354), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(KEYINPUT88), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT89), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n336), .A2(new_n351), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n336), .A2(new_n351), .A3(KEYINPUT75), .ZN(new_n530));
  AOI21_X1  g344(.A(G146), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT88), .B1(new_n531), .B2(new_n522), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n533));
  INV_X1    g347(.A(new_n525), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n513), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n517), .A2(KEYINPUT18), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n526), .A2(new_n535), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n505), .B(new_n520), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT19), .B1(new_n529), .B2(new_n530), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(KEYINPUT19), .B2(new_n527), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n191), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n548), .A2(new_n338), .A3(new_n514), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n526), .A2(new_n535), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT92), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n541), .A4(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n545), .B1(new_n554), .B2(new_n505), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n555), .A2(KEYINPUT20), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT20), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G122), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n560), .B2(G116), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n240), .B2(G122), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n560), .A2(KEYINPUT14), .A3(G116), .ZN(new_n563));
  OAI21_X1  g377(.A(G107), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT96), .ZN(new_n565));
  XNOR2_X1  g379(.A(G116), .B(G122), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n226), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT94), .B1(new_n202), .B2(G143), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n193), .A3(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n202), .A2(G143), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n571), .A2(new_n374), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n374), .B1(new_n571), .B2(new_n572), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n567), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT13), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n572), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n573), .B1(new_n584), .B2(G134), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n566), .B(new_n226), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n498), .A2(G217), .A3(new_n213), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n577), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n577), .B2(new_n587), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n291), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n552), .A2(new_n553), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n505), .B1(new_n597), .B2(new_n520), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n504), .B(new_n519), .C1(new_n552), .C2(new_n553), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n291), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G475), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n559), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(KEYINPUT97), .A2(G952), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(KEYINPUT97), .A2(G952), .ZN(new_n605));
  AOI21_X1  g419(.A(G953), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(G234), .A2(G237), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT21), .B(G898), .Z(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(G902), .A3(G953), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT98), .B1(new_n602), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n549), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n505), .B1(new_n597), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n556), .B1(new_n615), .B2(new_n599), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT20), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n555), .A2(KEYINPUT20), .A3(new_n556), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n601), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n611), .A4(new_n596), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n501), .B1(new_n613), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n316), .A2(new_n462), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND3_X1  g440(.A1(new_n308), .A2(new_n298), .A3(new_n309), .ZN(new_n627));
  INV_X1    g441(.A(new_n189), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n187), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n299), .A2(new_n311), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  OR3_X1    g448(.A1(new_n590), .A2(new_n591), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n634), .B1(new_n590), .B2(new_n591), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(G478), .A3(new_n291), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n592), .A2(new_n593), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n620), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n434), .A2(new_n291), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n436), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n644), .A2(new_n371), .A3(new_n501), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n633), .A2(new_n611), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND4_X1  g462(.A1(new_n601), .A2(new_n618), .A3(new_n595), .A4(new_n619), .ZN(new_n649));
  OR3_X1    g463(.A1(new_n649), .A2(KEYINPUT100), .A3(new_n612), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT100), .B1(new_n649), .B2(new_n612), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n633), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT35), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n226), .ZN(G9));
  INV_X1    g469(.A(new_n644), .ZN(new_n656));
  INV_X1    g470(.A(new_n369), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n348), .A2(new_n658), .A3(new_n355), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n658), .B1(new_n348), .B2(new_n355), .ZN(new_n661));
  OAI22_X1  g475(.A1(new_n660), .A2(new_n661), .B1(KEYINPUT36), .B2(new_n360), .ZN(new_n662));
  INV_X1    g476(.A(new_n661), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n659), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n657), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n367), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n316), .A2(new_n624), .A3(new_n656), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT102), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI21_X1  g486(.A(new_n501), .B1(new_n447), .B2(new_n461), .ZN(new_n673));
  INV_X1    g487(.A(new_n649), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n608), .B(KEYINPUT103), .Z(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(G900), .B2(new_n610), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n667), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n633), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  XOR2_X1   g495(.A(new_n677), .B(KEYINPUT39), .Z(new_n682));
  NOR2_X1   g496(.A1(new_n501), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n684), .B1(new_n501), .B2(new_n682), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n187), .A3(new_n687), .A4(new_n667), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n627), .A2(new_n628), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n690), .A2(KEYINPUT38), .A3(new_n310), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT38), .B1(new_n690), .B2(new_n310), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n620), .A2(new_n595), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n445), .A2(new_n446), .ZN(new_n696));
  INV_X1    g510(.A(G472), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n404), .A2(new_n410), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n455), .B2(new_n410), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n697), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n440), .A2(new_n441), .ZN(new_n703));
  AOI211_X1 g517(.A(KEYINPUT69), .B(KEYINPUT32), .C1(new_n434), .C2(new_n435), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n696), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n689), .A2(new_n693), .A3(new_n695), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  AND3_X1   g521(.A1(new_n620), .A2(new_n639), .A3(new_n677), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n633), .A2(new_n668), .A3(new_n673), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  OAI211_X1 g524(.A(new_n696), .B(new_n461), .C1(new_n703), .C2(new_n704), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n291), .B1(new_n487), .B2(new_n491), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n463), .A2(KEYINPUT105), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n714), .A2(new_n500), .A3(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n711), .A2(new_n370), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n633), .A3(new_n611), .A4(new_n641), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT41), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G113), .ZN(G15));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n633), .A3(new_n652), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND2_X1  g536(.A1(new_n613), .A2(new_n623), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n667), .B1(new_n447), .B2(new_n461), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n633), .A2(new_n723), .A3(new_n716), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI21_X1  g540(.A(new_n415), .B1(new_n411), .B2(new_n457), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n435), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n642), .B2(G472), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n730), .B(new_n697), .C1(new_n434), .C2(new_n291), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n370), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n716), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(new_n694), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n633), .A2(new_n611), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  OAI211_X1 g550(.A(new_n668), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n620), .A2(new_n639), .A3(new_n677), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n633), .A2(new_n716), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(new_n501), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n690), .A2(new_n310), .A3(new_n187), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n711), .A3(new_n370), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n690), .A2(new_n310), .A3(new_n187), .A4(new_n742), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n461), .A2(new_n438), .A3(new_n443), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n370), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n746), .A2(new_n748), .A3(new_n738), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT42), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n381), .ZN(G33));
  NAND2_X1  g566(.A1(new_n711), .A2(new_n370), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n678), .A3(new_n746), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n374), .ZN(G36));
  NAND4_X1  g569(.A1(new_n559), .A2(KEYINPUT43), .A3(new_n601), .A4(new_n639), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n601), .A2(new_n618), .A3(new_n639), .A4(new_n619), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n644), .A3(new_n668), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n690), .A2(new_n310), .A3(new_n187), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n760), .A2(KEYINPUT44), .A3(new_n644), .A4(new_n668), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  INV_X1    g582(.A(new_n486), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT78), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n234), .B2(new_n387), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n469), .A3(new_n480), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT12), .B1(new_n772), .B2(new_n383), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n489), .B1(new_n769), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n468), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT45), .B1(new_n775), .B2(new_n494), .ZN(new_n776));
  OAI211_X1 g590(.A(KEYINPUT45), .B(new_n494), .C1(new_n495), .C2(new_n488), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n768), .B(G469), .C1(new_n779), .C2(G902), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n496), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(G469), .A3(new_n777), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n493), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n492), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n682), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n500), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n767), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(new_n500), .ZN(new_n790));
  INV_X1    g604(.A(new_n492), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n783), .A2(new_n493), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n791), .B1(new_n792), .B2(new_n768), .ZN(new_n793));
  AOI211_X1 g607(.A(KEYINPUT47), .B(new_n790), .C1(new_n793), .C2(new_n784), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n785), .B2(new_n500), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n764), .A2(new_n738), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n711), .A2(new_n370), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n718), .A2(new_n725), .A3(new_n721), .A4(new_n735), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n559), .A2(new_n805), .A3(new_n595), .A4(new_n601), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n649), .A2(KEYINPUT108), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n807), .A3(new_n640), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n808), .A2(new_n645), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n316), .A2(new_n611), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n625), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n677), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n620), .A2(new_n595), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n711), .A2(new_n668), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n643), .A2(new_n730), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n642), .A2(KEYINPUT106), .A3(G472), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n708), .A2(new_n668), .A3(new_n728), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n746), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n751), .A2(new_n754), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n804), .A2(new_n811), .A3(new_n820), .A4(new_n669), .ZN(new_n821));
  INV_X1    g635(.A(new_n187), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n299), .B2(KEYINPUT99), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n690), .A2(new_n632), .A3(new_n310), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n711), .A2(new_n823), .A3(new_n742), .A4(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n716), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n825), .A2(new_n679), .B1(new_n826), .B2(new_n739), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT109), .B1(new_n667), .B2(new_n677), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT109), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n367), .A2(new_n666), .A3(new_n830), .A4(new_n812), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n742), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n447), .B2(new_n702), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n824), .A3(new_n823), .A4(new_n695), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n827), .A2(new_n828), .A3(new_n709), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n709), .A2(new_n680), .A3(new_n740), .A4(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n802), .B1(new_n821), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n669), .A2(new_n625), .A3(new_n810), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n814), .A2(new_n818), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n743), .ZN(new_n843));
  INV_X1    g657(.A(new_n748), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n743), .A2(new_n708), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT42), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n462), .A2(new_n674), .A3(new_n677), .A4(new_n743), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n846), .A3(new_n745), .A4(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n841), .A2(new_n803), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n837), .A4(new_n835), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n839), .A2(new_n840), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n840), .B1(new_n839), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n760), .A2(new_n675), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n690), .A2(new_n310), .A3(new_n716), .A4(new_n187), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n737), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n676), .B1(new_n756), .B2(new_n759), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n732), .A2(new_n733), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n859), .A2(new_n860), .A3(new_n822), .ZN(new_n861));
  INV_X1    g675(.A(new_n693), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT50), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n859), .A2(new_n860), .A3(new_n822), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n693), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n858), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n856), .A2(new_n705), .ZN(new_n868));
  INV_X1    g682(.A(new_n608), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n370), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT110), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n856), .A2(new_n705), .A3(new_n873), .A4(new_n870), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n620), .A2(new_n639), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT111), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT110), .B1(new_n868), .B2(new_n871), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n875), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(KEYINPUT111), .A3(new_n877), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n867), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n855), .A2(new_n732), .A3(new_n764), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n714), .A2(new_n715), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n790), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n794), .B2(new_n796), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT51), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(KEYINPUT112), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n887), .B(new_n892), .C1(new_n794), .C2(new_n796), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n885), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(KEYINPUT51), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT50), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n865), .B1(new_n864), .B2(new_n693), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n857), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(KEYINPUT111), .A2(new_n874), .A3(new_n876), .A4(new_n877), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT111), .B1(new_n882), .B2(new_n877), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n882), .A2(new_n641), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n633), .A2(new_n860), .A3(new_n859), .ZN(new_n903));
  INV_X1    g717(.A(new_n606), .ZN(new_n904));
  INV_X1    g718(.A(new_n856), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n859), .A3(new_n844), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT48), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n859), .A3(new_n908), .A4(new_n844), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT113), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n889), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT113), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n901), .A4(new_n912), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n853), .A2(new_n854), .A3(new_n914), .A4(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n821), .A2(new_n838), .A3(new_n802), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n836), .B(new_n828), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n922), .B2(new_n849), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n839), .A2(new_n850), .A3(new_n840), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n924), .A2(new_n914), .A3(new_n925), .A4(new_n919), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT114), .ZN(new_n927));
  OR2_X1    g741(.A1(G952), .A2(G953), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n920), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n886), .B(KEYINPUT49), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n705), .ZN(new_n931));
  INV_X1    g745(.A(new_n757), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n370), .A2(new_n188), .A3(new_n500), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT107), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n862), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n213), .A2(G952), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(G210), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n939), .B(new_n291), .C1(new_n839), .C2(new_n850), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(KEYINPUT56), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n296), .B(KEYINPUT115), .Z(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(new_n297), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n938), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT117), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n940), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n839), .A2(new_n850), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(new_n948), .A3(G210), .A4(G902), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n945), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT118), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(G210), .B(G902), .C1(new_n921), .C2(new_n923), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT56), .B1(new_n954), .B2(KEYINPUT117), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT118), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n956), .A3(new_n951), .A4(new_n945), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n946), .B1(new_n953), .B2(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n493), .B(KEYINPUT57), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n853), .A2(new_n959), .B1(new_n491), .B2(new_n487), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n783), .B(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n950), .A2(G902), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n937), .B1(new_n960), .B2(new_n962), .ZN(G54));
  INV_X1    g777(.A(KEYINPUT58), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n964), .B(new_n291), .C1(new_n839), .C2(new_n850), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n555), .B1(new_n965), .B2(G475), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n968));
  INV_X1    g782(.A(new_n555), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n965), .A2(KEYINPUT120), .A3(G475), .A4(new_n555), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n937), .B(new_n966), .C1(new_n970), .C2(new_n971), .ZN(G60));
  NAND2_X1  g786(.A1(new_n635), .A2(new_n636), .ZN(new_n973));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT59), .Z(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n853), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n977), .B(new_n978), .C1(new_n851), .C2(new_n852), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n976), .A2(new_n938), .A3(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  NAND2_X1  g796(.A1(new_n950), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n368), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n937), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n662), .A2(new_n665), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n983), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n985), .B(KEYINPUT61), .C1(new_n986), .C2(new_n983), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(G66));
  NAND3_X1  g805(.A1(new_n609), .A2(G953), .A3(new_n212), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n841), .A2(new_n803), .A3(KEYINPUT121), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT121), .B1(new_n841), .B2(new_n803), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n995), .B2(G953), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n942), .B1(G898), .B2(new_n213), .ZN(new_n997));
  XOR2_X1   g811(.A(KEYINPUT122), .B(KEYINPUT123), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n996), .B(new_n999), .ZN(G69));
  INV_X1    g814(.A(G900), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n464), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n403), .B(new_n547), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n213), .A2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n633), .A2(new_n695), .A3(new_n844), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n787), .B1(new_n767), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n709), .A2(new_n680), .A3(new_n740), .A4(new_n847), .ZN(new_n1009));
  INV_X1    g823(.A(new_n800), .ZN(new_n1010));
  NOR4_X1   g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n751), .A4(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1006), .B1(new_n1011), .B2(G953), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT125), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT125), .B(new_n1006), .C1(new_n1011), .C2(G953), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1002), .B1(new_n1016), .B2(KEYINPUT124), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n462), .A2(new_n683), .A3(new_n765), .A4(new_n808), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n788), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n827), .A2(new_n706), .A3(new_n709), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n1019), .B(new_n800), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1003), .B1(new_n1024), .B2(new_n213), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1017), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1028));
  AOI221_X4 g842(.A(new_n1025), .B1(KEYINPUT124), .B2(new_n1002), .C1(new_n1028), .C2(new_n1003), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1027), .A2(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  INV_X1    g846(.A(new_n451), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n450), .A2(new_n410), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT127), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1036), .B1(new_n839), .B2(new_n850), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n1024), .A2(new_n995), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n699), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n993), .A2(new_n1011), .A3(new_n994), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1032), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1041), .A2(new_n404), .A3(new_n410), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(new_n938), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(KEYINPUT126), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT126), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1042), .A2(new_n1045), .A3(new_n938), .ZN(new_n1046));
  AOI211_X1 g860(.A(new_n1037), .B(new_n1039), .C1(new_n1044), .C2(new_n1046), .ZN(G57));
endmodule


