//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1386, new_n1387;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n208), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n217), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n225), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n226), .A2(G33), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n251), .A2(new_n202), .B1(new_n226), .B2(G68), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n226), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G50), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n250), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT11), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n250), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G1), .B2(new_n226), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT12), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n262), .B1(new_n265), .B2(new_n210), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n264), .A2(KEYINPUT12), .A3(G68), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n261), .A2(new_n210), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n257), .A2(new_n258), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n259), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(G274), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT67), .B(G45), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G41), .A2(G45), .ZN(new_n279));
  OAI22_X1  g0079(.A1(new_n278), .A2(new_n225), .B1(new_n279), .B2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n277), .B1(new_n287), .B2(G238), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(G232), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  OAI211_X1 g0092(.A(G226), .B(new_n292), .C1(new_n289), .C2(new_n290), .ZN(new_n293));
  AND3_X1   g0093(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT72), .B1(G33), .B2(G97), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n278), .A2(new_n225), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n272), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n284), .B1(new_n283), .B2(new_n285), .ZN(new_n302));
  OAI21_X1  g0102(.A(G238), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n299), .A2(new_n303), .A3(new_n272), .A4(new_n276), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n300), .A2(new_n305), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(KEYINPUT14), .B1(new_n307), .B2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n303), .A3(new_n276), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  AOI211_X1 g0111(.A(KEYINPUT14), .B(new_n309), .C1(new_n311), .C2(new_n304), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT73), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(G179), .A3(new_n304), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n309), .B1(new_n311), .B2(new_n304), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(new_n312), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n271), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n271), .B1(new_n307), .B2(G190), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n307), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n277), .B1(new_n287), .B2(G226), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n253), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n292), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n289), .A2(new_n290), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(G223), .B1(new_n331), .B2(G77), .ZN(new_n332));
  AOI21_X1  g0132(.A(G1698), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G222), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n326), .B1(new_n335), .B2(new_n283), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n336), .A2(G200), .B1(KEYINPUT71), .B2(KEYINPUT10), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n251), .ZN(new_n341));
  INV_X1    g0141(.A(G150), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n201), .A2(new_n226), .B1(new_n254), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n250), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n265), .A2(new_n255), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(new_n255), .C2(new_n261), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT9), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n338), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT10), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n348), .B(new_n351), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n336), .A2(G179), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n336), .A2(new_n309), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g0156(.A(G232), .B(new_n292), .C1(new_n289), .C2(new_n290), .ZN(new_n357));
  OAI211_X1 g0157(.A(G238), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n328), .A2(G107), .A3(new_n329), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n298), .ZN(new_n361));
  OAI21_X1  g0161(.A(G244), .B1(new_n301), .B2(new_n302), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(new_n276), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT69), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT69), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(new_n276), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(G200), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G20), .A2(G77), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT15), .B(G87), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n340), .B2(new_n254), .C1(new_n251), .C2(new_n369), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n370), .A2(new_n250), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n265), .A2(new_n202), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n261), .B2(new_n202), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n277), .B1(new_n287), .B2(G244), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n365), .B1(new_n376), .B2(new_n361), .ZN(new_n377));
  AND4_X1   g0177(.A1(new_n365), .A2(new_n361), .A3(new_n276), .A4(new_n362), .ZN(new_n378));
  OAI21_X1  g0178(.A(G190), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT70), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n364), .A2(new_n366), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(G190), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n375), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n374), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n364), .A2(new_n309), .A3(new_n366), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n325), .A2(new_n356), .A3(new_n384), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n328), .A2(new_n226), .A3(new_n329), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n328), .A2(new_n394), .A3(new_n226), .A4(new_n329), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(G68), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT76), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(G68), .A4(new_n395), .ZN(new_n399));
  XNOR2_X1  g0199(.A(G58), .B(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G20), .A2(G33), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n400), .A2(G20), .B1(G159), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n396), .A2(KEYINPUT74), .A3(KEYINPUT16), .A4(new_n402), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n410), .A3(new_n250), .ZN(new_n411));
  INV_X1    g0211(.A(new_n340), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n265), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n412), .B2(new_n261), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(G226), .B2(new_n292), .C1(new_n289), .C2(new_n290), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n283), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(G190), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n280), .A2(new_n217), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT77), .B1(new_n277), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT77), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(new_n276), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(new_n276), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n323), .B1(new_n427), .B2(new_n419), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AND4_X1   g0229(.A1(KEYINPUT17), .A2(new_n411), .A3(new_n415), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n260), .B1(new_n408), .B2(new_n409), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n414), .B1(new_n431), .B2(new_n405), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT17), .B1(new_n432), .B2(new_n429), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n391), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n411), .A2(new_n415), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n419), .A2(G179), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n422), .A3(new_n425), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n309), .B1(new_n427), .B2(new_n419), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n432), .A2(new_n440), .A3(KEYINPUT18), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n411), .A2(new_n415), .A3(new_n429), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT17), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(KEYINPUT78), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n434), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n390), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n292), .B1(new_n289), .B2(new_n290), .ZN(new_n454));
  OAI21_X1  g0254(.A(G244), .B1(KEYINPUT81), .B2(KEYINPUT4), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n328), .A2(new_n329), .ZN(new_n457));
  INV_X1    g0257(.A(new_n455), .ZN(new_n458));
  INV_X1    g0258(.A(new_n453), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n457), .A2(new_n292), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n330), .A2(G250), .ZN(new_n461));
  NAND3_X1  g0261(.A1(KEYINPUT82), .A2(G33), .A3(G283), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT82), .B1(G33), .B2(G283), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n456), .A2(new_n460), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(G250), .B2(new_n330), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT83), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n460), .A4(new_n456), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n471), .A3(new_n298), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n298), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G257), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(G274), .A3(new_n283), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(G190), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n283), .B1(new_n467), .B2(KEYINPUT83), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n479), .B1(new_n484), .B2(new_n471), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .A3(G190), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n323), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n264), .A2(G97), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n264), .B1(G1), .B2(new_n253), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(new_n250), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(G97), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n393), .A2(G107), .A3(new_n395), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  AND2_X1   g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G20), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n401), .A2(G77), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT79), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n493), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT80), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n250), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n505), .B2(new_n250), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n492), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n488), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n492), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n505), .A2(new_n250), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(new_n507), .ZN(new_n515));
  AOI21_X1  g0315(.A(G169), .B1(new_n472), .B2(new_n480), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n485), .A2(new_n385), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n487), .A2(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n264), .A2(G116), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n491), .B2(G116), .ZN(new_n522));
  AOI21_X1  g0322(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n463), .B2(new_n464), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n249), .A2(new_n225), .B1(G20), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT20), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n475), .A2(new_n474), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G270), .A3(new_n283), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n478), .ZN(new_n533));
  OAI211_X1 g0333(.A(G264), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n328), .A2(G303), .A3(new_n329), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(new_n454), .C2(new_n219), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n283), .B1(new_n536), .B2(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n333), .A2(G257), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT88), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n534), .A4(new_n535), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n520), .B1(new_n530), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(KEYINPUT88), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n298), .A3(new_n540), .ZN(new_n544));
  INV_X1    g0344(.A(new_n533), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n524), .A2(new_n526), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n526), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n309), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n552), .A3(KEYINPUT21), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n541), .A2(G179), .A3(new_n529), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n542), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n529), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n541), .B2(new_n323), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n337), .B(new_n533), .C1(new_n537), .C2(new_n540), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n474), .B(KEYINPUT85), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n298), .A2(new_n213), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(G45), .B2(new_n274), .ZN(new_n563));
  OAI211_X1 g0363(.A(G244), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT86), .B1(new_n454), .B2(new_n211), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT86), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n333), .A2(new_n568), .A3(G238), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n563), .B1(new_n570), .B2(new_n283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT72), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G87), .A2(G97), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n579), .A2(KEYINPUT87), .A3(new_n498), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT87), .B1(new_n579), .B2(new_n498), .ZN(new_n581));
  OAI22_X1  g0381(.A1(new_n578), .A2(G20), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n226), .B(G68), .C1(new_n289), .C2(new_n290), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n251), .B2(new_n218), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n260), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n490), .A2(new_n212), .A3(new_n250), .ZN(new_n587));
  INV_X1    g0387(.A(new_n369), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n588), .A2(new_n264), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G190), .B(new_n563), .C1(new_n570), .C2(new_n283), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n572), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n571), .A2(new_n309), .ZN(new_n593));
  INV_X1    g0393(.A(new_n589), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n491), .A2(new_n588), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n582), .A2(new_n585), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n260), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n385), .B(new_n563), .C1(new_n570), .C2(new_n283), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n226), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT22), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n457), .A2(new_n603), .A3(new_n226), .A4(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT24), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n565), .A2(G20), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n226), .B2(G107), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n498), .A2(KEYINPUT23), .A3(G20), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n605), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n250), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g0414(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n615));
  NOR2_X1   g0415(.A1(new_n264), .A2(G107), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(G107), .B2(new_n491), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT90), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(G294), .ZN(new_n621));
  INV_X1    g0421(.A(G294), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(KEYINPUT90), .ZN(new_n623));
  OAI21_X1  g0423(.A(G33), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(G250), .B(new_n292), .C1(new_n289), .C2(new_n290), .ZN(new_n625));
  OAI211_X1 g0425(.A(G257), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n298), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n476), .A2(G264), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n478), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(G190), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n627), .A2(new_n298), .B1(new_n476), .B2(G264), .ZN(new_n632));
  AOI21_X1  g0432(.A(G200), .B1(new_n632), .B2(new_n478), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT91), .B1(new_n619), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n323), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(G190), .B2(new_n630), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT91), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n614), .A4(new_n618), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n600), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n309), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n632), .A2(new_n385), .A3(new_n478), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n619), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n519), .A2(new_n560), .A3(new_n640), .A4(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n452), .A2(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n452), .ZN(new_n646));
  INV_X1    g0446(.A(new_n599), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n592), .A2(new_n599), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n517), .A4(new_n518), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n472), .A2(new_n480), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n309), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n518), .A3(new_n510), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n653), .B2(new_n600), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n647), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n487), .A2(new_n511), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n643), .A2(new_n542), .A3(new_n553), .A4(new_n554), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n640), .A2(new_n656), .A3(new_n653), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n355), .ZN(new_n661));
  INV_X1    g0461(.A(new_n321), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n389), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n434), .A2(new_n449), .A3(new_n324), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n444), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n661), .B1(new_n665), .B2(new_n352), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n263), .A2(new_n226), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G343), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n529), .ZN(new_n674));
  MUX2_X1   g0474(.A(new_n555), .B(new_n560), .S(new_n674), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n635), .A2(new_n639), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n614), .B2(new_n618), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n643), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n643), .A2(new_n673), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n680), .A2(new_n555), .A3(new_n643), .A4(new_n672), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0488(.A(new_n229), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n580), .A2(new_n581), .A3(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(G1), .ZN(new_n693));
  INV_X1    g0493(.A(new_n224), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n691), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n658), .A2(KEYINPUT96), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT95), .ZN(new_n698));
  NOR4_X1   g0498(.A1(new_n653), .A2(new_n600), .A3(new_n698), .A4(new_n650), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n647), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n649), .A2(new_n654), .A3(new_n698), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n519), .A2(new_n702), .A3(new_n640), .A4(new_n657), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n697), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n672), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n659), .A2(new_n672), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n677), .A2(new_n560), .A3(new_n648), .A4(new_n643), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n656), .A2(new_n653), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n713), .A3(new_n673), .ZN(new_n714));
  INV_X1    g0514(.A(new_n632), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n571), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n385), .B(new_n533), .C1(new_n537), .C2(new_n540), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n485), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n485), .A2(new_n716), .A3(new_n717), .A4(KEYINPUT30), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n632), .B2(new_n478), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n546), .A2(new_n723), .A3(new_n571), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n722), .B1(new_n724), .B2(new_n485), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n571), .A2(new_n385), .A3(new_n630), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n651), .A3(KEYINPUT93), .A4(new_n546), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n720), .A2(new_n721), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n673), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(new_n651), .A3(new_n546), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n720), .A2(new_n721), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n672), .A2(new_n730), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n714), .B1(new_n736), .B2(KEYINPUT94), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT94), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n731), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n711), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n710), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n696), .B1(new_n743), .B2(G1), .ZN(G364));
  NAND2_X1  g0544(.A1(new_n226), .A2(G13), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n263), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n690), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n675), .B2(G330), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G330), .B2(new_n675), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n689), .A2(new_n331), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n753), .A2(new_n206), .B1(G116), .B2(new_n229), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n689), .A2(new_n457), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n247), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n275), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n224), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n754), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n225), .B1(G20), .B2(new_n309), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  OAI21_X1  g0566(.A(new_n749), .B1(new_n760), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n226), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n226), .A2(new_n337), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n385), .A2(new_n323), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n323), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n768), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n777), .A2(G50), .B1(new_n780), .B2(G107), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n774), .A2(new_n778), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n773), .B(new_n781), .C1(new_n212), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n226), .B1(new_n769), .B2(G190), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n218), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n385), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n457), .B1(new_n787), .B2(new_n216), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(new_n768), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n768), .A2(new_n786), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n210), .B1(new_n790), .B2(new_n202), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n783), .A2(new_n785), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT98), .Z(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n794), .A2(new_n789), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n787), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n457), .B(new_n796), .C1(G322), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n621), .A2(new_n623), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n784), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(new_n777), .B2(G326), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  INV_X1    g0605(.A(G329), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n779), .A2(new_n805), .B1(new_n770), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n782), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(G303), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n798), .A2(new_n803), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n793), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n767), .B1(new_n811), .B2(new_n764), .ZN(new_n812));
  INV_X1    g0612(.A(new_n763), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n675), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n751), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  INV_X1    g0616(.A(KEYINPUT101), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n374), .A2(new_n672), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n384), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n673), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n817), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n367), .A2(new_n374), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n382), .B1(new_n381), .B2(G190), .ZN(new_n825));
  AOI211_X1 g0625(.A(KEYINPUT70), .B(new_n337), .C1(new_n364), .C2(new_n366), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n819), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n389), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n829), .A2(KEYINPUT101), .A3(new_n821), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n707), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT101), .B1(new_n829), .B2(new_n821), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n820), .A2(new_n817), .A3(new_n822), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n659), .A2(new_n672), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n740), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT102), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n740), .B1(new_n831), .B2(new_n834), .ZN(new_n839));
  OR4_X1    g0639(.A1(new_n749), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n749), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n764), .A2(new_n761), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n202), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n764), .ZN(new_n844));
  INV_X1    g0644(.A(new_n789), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G283), .A2(new_n845), .B1(new_n846), .B2(G116), .ZN(new_n847));
  INV_X1    g0647(.A(G303), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n776), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT100), .Z(new_n850));
  AOI22_X1  g0650(.A1(G107), .A2(new_n808), .B1(new_n797), .B2(G294), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n795), .B2(new_n770), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n331), .B1(new_n779), .B2(new_n212), .ZN(new_n853));
  NOR4_X1   g0653(.A1(new_n850), .A2(new_n785), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G137), .A2(new_n777), .B1(new_n845), .B2(G150), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n797), .B1(new_n846), .B2(G159), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n457), .B1(new_n782), .B2(new_n255), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n779), .A2(new_n210), .B1(new_n770), .B2(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n859), .B(new_n861), .C1(G58), .C2(new_n801), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n857), .A2(KEYINPUT34), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n854), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n830), .A2(new_n823), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n843), .B1(new_n844), .B2(new_n866), .C1(new_n867), .C2(new_n762), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n840), .A2(new_n868), .ZN(G384));
  OR2_X1    g0669(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(G116), .A4(new_n227), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  OAI211_X1 g0673(.A(new_n224), .B(G77), .C1(new_n216), .C2(new_n210), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n255), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n263), .B(G13), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AOI221_X4 g0677(.A(new_n414), .B1(new_n428), .B2(new_n426), .C1(new_n431), .C2(new_n405), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n671), .B1(new_n438), .B2(new_n439), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n411), .B2(new_n415), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT107), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT107), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n445), .B(new_n882), .C1(new_n432), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT106), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n436), .A2(new_n435), .A3(new_n441), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT18), .B1(new_n432), .B2(new_n440), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n890), .A2(new_n447), .A3(new_n891), .A4(new_n448), .ZN(new_n892));
  INV_X1    g0692(.A(new_n671), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n432), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n888), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n881), .A3(new_n883), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n889), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n396), .A2(new_n402), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n404), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n414), .B1(new_n431), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n893), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n450), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n445), .B1(new_n903), .B2(new_n879), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT103), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n909), .A3(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(new_n880), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n445), .A3(new_n885), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n905), .A2(new_n913), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n899), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n662), .A2(new_n672), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n834), .A2(new_n822), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n270), .A2(new_n672), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n321), .A2(new_n324), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n314), .B2(new_n320), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n905), .B2(new_n913), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT105), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n919), .A2(new_n934), .A3(new_n914), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n930), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n444), .A2(new_n671), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n923), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n709), .A2(new_n646), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n666), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n938), .B(new_n940), .Z(new_n941));
  NAND3_X1  g0741(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n731), .B(new_n942), .C1(new_n644), .C2(new_n673), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n929), .A2(new_n867), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT105), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n934), .B1(new_n919), .B2(new_n914), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n900), .A2(new_n914), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n929), .A2(new_n867), .A3(new_n943), .A4(KEYINPUT40), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT108), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g0751(.A1(KEYINPUT40), .A2(new_n929), .A3(new_n867), .A4(new_n943), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT108), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n953), .A3(new_n915), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n947), .A2(new_n948), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n640), .A2(new_n643), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n956), .A2(new_n519), .A3(new_n560), .A4(new_n672), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n731), .A2(new_n942), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n452), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n711), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n959), .B2(new_n955), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n941), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n263), .B2(new_n746), .C1(new_n941), .C2(new_n961), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n962), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n877), .B1(new_n965), .B2(new_n966), .ZN(G367));
  OAI21_X1  g0767(.A(new_n519), .B1(new_n515), .B2(new_n672), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT110), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(KEYINPUT110), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n653), .B1(new_n971), .B2(new_n643), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n672), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n517), .A2(new_n518), .A3(new_n673), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n974), .A3(new_n970), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT42), .B1(new_n976), .B2(new_n685), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT42), .ZN(new_n978));
  INV_X1    g0778(.A(new_n685), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n590), .A2(new_n672), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n600), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n647), .A2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT43), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n981), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n977), .A2(new_n980), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n991), .A2(new_n987), .A3(new_n986), .A4(new_n973), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n976), .A2(new_n684), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n990), .B2(new_n992), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n690), .B(KEYINPUT41), .Z(new_n997));
  AND3_X1   g0797(.A1(new_n975), .A2(KEYINPUT45), .A3(new_n686), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT45), .B1(new_n975), .B2(new_n686), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT111), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1001), .B(KEYINPUT44), .C1(new_n975), .C2(new_n686), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n686), .B1(KEYINPUT111), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(KEYINPUT44), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n976), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1000), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n683), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1000), .A2(new_n684), .A3(new_n1002), .A4(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n555), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n682), .B1(new_n1010), .B2(new_n673), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n685), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n676), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n742), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1008), .A2(new_n1009), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n997), .B1(new_n1015), .B2(new_n743), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n996), .B1(new_n1016), .B2(new_n748), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n766), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n229), .B2(new_n369), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n240), .A2(new_n756), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n749), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n808), .A2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n800), .A2(new_n845), .B1(new_n797), .B2(G303), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n805), .C2(new_n790), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n779), .A2(new_n218), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G311), .B2(new_n777), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n770), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n457), .B1(new_n1028), .B2(G317), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(new_n498), .C2(new_n784), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n779), .A2(new_n202), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G137), .B2(new_n1028), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n255), .B2(new_n790), .C1(new_n771), .C2(new_n789), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G143), .A2(new_n777), .B1(new_n808), .B2(G58), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n801), .A2(G68), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n331), .B1(new_n797), .B2(G150), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1025), .A2(new_n1030), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1021), .B1(new_n1039), .B2(new_n764), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n813), .B2(new_n985), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1017), .A2(new_n1041), .ZN(G387));
  NOR2_X1   g0842(.A1(new_n1013), .A2(new_n747), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n753), .A2(new_n692), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n237), .A2(new_n758), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n755), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n692), .B(new_n473), .C1(new_n210), .C2(new_n202), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT50), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n340), .B2(G50), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n412), .A2(KEYINPUT50), .A3(new_n255), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1046), .A2(new_n1051), .B1(G107), .B2(new_n229), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n841), .B1(new_n1052), .B2(new_n1018), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n457), .B1(new_n1028), .B2(G326), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n799), .A2(new_n782), .B1(new_n784), .B2(new_n805), .ZN(new_n1055));
  INV_X1    g0855(.A(G322), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n776), .A2(new_n1056), .B1(new_n789), .B2(new_n795), .ZN(new_n1057));
  INV_X1    g0857(.A(G317), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n787), .A2(new_n1058), .B1(new_n790), .B2(new_n848), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1055), .B1(new_n1060), .B2(KEYINPUT48), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT48), .B2(new_n1060), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1054), .B1(new_n525), .B2(new_n779), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n784), .A2(new_n369), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G50), .B2(new_n797), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT112), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G68), .A2(new_n846), .B1(new_n1028), .B2(G150), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n340), .B2(new_n789), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n776), .A2(new_n771), .B1(new_n782), .B2(new_n202), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1070), .A2(new_n331), .A3(new_n1026), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1065), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1053), .B1(new_n1073), .B2(new_n844), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n682), .B2(new_n763), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1043), .A2(new_n1075), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n742), .A2(new_n1013), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n690), .B1(new_n742), .B2(new_n1013), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n1008), .A2(new_n748), .A3(new_n1009), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1018), .B1(new_n218), .B2(new_n229), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n244), .A2(new_n755), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n749), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n782), .A2(new_n805), .B1(new_n770), .B2(new_n1056), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT113), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n331), .B1(new_n779), .B2(new_n498), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n789), .A2(new_n848), .B1(new_n790), .B2(new_n622), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G116), .C2(new_n801), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n776), .A2(new_n1058), .B1(new_n787), .B2(new_n795), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n776), .A2(new_n342), .B1(new_n787), .B2(new_n771), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n845), .A2(G50), .B1(new_n846), .B2(new_n412), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G68), .A2(new_n808), .B1(new_n1028), .B2(G143), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n784), .A2(new_n202), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n331), .B(new_n1099), .C1(G87), .C2(new_n780), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1083), .B1(new_n1102), .B2(new_n764), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n975), .B2(new_n813), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1015), .A2(new_n690), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1014), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1080), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(G390));
  AOI21_X1  g0907(.A(KEYINPUT31), .B1(new_n728), .B2(new_n673), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n733), .A2(new_n734), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT94), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n739), .A2(new_n1110), .A3(new_n957), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(G330), .A3(new_n867), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT116), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n929), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n944), .A2(G330), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1113), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n924), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n711), .B1(new_n958), .B2(new_n957), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n929), .B1(new_n1120), .B2(new_n867), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n704), .A2(new_n867), .A3(new_n672), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n822), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1111), .A2(G330), .A3(new_n867), .A4(new_n929), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT115), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1119), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n740), .A2(KEYINPUT115), .A3(new_n867), .A4(new_n929), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1127), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1123), .A2(new_n929), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n915), .A2(new_n922), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n673), .B1(new_n655), .B2(new_n658), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n821), .B1(new_n867), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n922), .B1(new_n1138), .B2(new_n1114), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n931), .A2(new_n932), .A3(new_n916), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT39), .B1(new_n900), .B2(new_n914), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1133), .A2(new_n1136), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1116), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n917), .A2(new_n920), .B1(new_n930), .B2(new_n922), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1114), .B1(new_n1122), .B2(new_n822), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n915), .A2(new_n922), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n646), .A2(new_n1120), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n939), .A2(new_n666), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1131), .A2(new_n1143), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n690), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT117), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1149), .A2(new_n1143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT116), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1116), .A3(new_n1115), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1160), .A2(new_n924), .B1(new_n1133), .B2(new_n1124), .ZN(new_n1161));
  OAI21_X1  g0961(.A(KEYINPUT118), .B1(new_n1161), .B2(new_n1151), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1151), .B1(new_n1119), .B2(new_n1130), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1157), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT117), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1153), .A2(new_n1167), .A3(new_n690), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1155), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1156), .A2(new_n748), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n921), .A2(new_n761), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n808), .A2(G150), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G159), .B2(new_n801), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  INV_X1    g0975(.A(G125), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n790), .A2(new_n1175), .B1(new_n770), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G50), .B2(new_n780), .ZN(new_n1178));
  INV_X1    g0978(.A(G137), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n860), .A2(new_n787), .B1(new_n789), .B2(new_n1179), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n331), .B(new_n1180), .C1(G128), .C2(new_n777), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n789), .A2(new_n498), .B1(new_n790), .B2(new_n218), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT119), .Z(new_n1184));
  AOI22_X1  g0984(.A1(G116), .A2(new_n797), .B1(new_n780), .B2(G68), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n777), .A2(G283), .B1(new_n1028), .B2(G294), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n457), .B(new_n1099), .C1(G87), .C2(new_n808), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n844), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n841), .B(new_n1189), .C1(new_n340), .C2(new_n842), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1171), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1170), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(G378));
  OAI22_X1  g0994(.A1(new_n776), .A2(new_n1176), .B1(new_n789), .B2(new_n860), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n846), .A2(G137), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n787), .C1(new_n782), .C2(new_n1175), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(G150), .C2(new_n801), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n779), .A2(new_n771), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G33), .A2(G41), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT120), .Z(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G124), .C2(new_n1028), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G116), .A2(new_n777), .B1(new_n808), .B2(G77), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n457), .A2(G41), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n780), .A2(G58), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n1035), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n218), .A2(new_n789), .B1(new_n787), .B2(new_n498), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n790), .A2(new_n369), .B1(new_n770), .B2(new_n805), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(KEYINPUT58), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1205), .B(new_n255), .C1(G41), .C2(new_n457), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1207), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n764), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n841), .B1(new_n255), .B2(new_n842), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n346), .A2(new_n671), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n356), .B(new_n1221), .Z(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1219), .B(new_n1220), .C1(new_n1225), .C2(new_n762), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n938), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1225), .B1(new_n955), .B2(G330), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n929), .A2(new_n867), .A3(new_n943), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n933), .B2(new_n935), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n949), .A2(KEYINPUT108), .A3(new_n950), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n953), .B1(new_n952), .B2(new_n915), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1231), .A2(KEYINPUT40), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1234), .A2(new_n711), .A3(new_n1224), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1224), .B1(new_n1234), .B2(new_n711), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n947), .A2(new_n948), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n951), .A2(new_n954), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1238), .A2(G330), .A3(new_n1239), .A4(new_n1225), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n938), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1227), .B1(new_n1242), .B2(new_n748), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1153), .A2(new_n1152), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1237), .A2(new_n938), .A3(new_n1240), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n938), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1246));
  OAI211_X1 g1046(.A(KEYINPUT57), .B(new_n1244), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n690), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1243), .B1(new_n1248), .B2(new_n1249), .ZN(G375));
  INV_X1    g1050(.A(new_n997), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1119), .A2(new_n1151), .A3(new_n1130), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1162), .A2(new_n1165), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n747), .B1(new_n1119), .B2(new_n1130), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n841), .B1(new_n210), .B2(new_n842), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n776), .A2(new_n860), .B1(new_n787), .B2(new_n1179), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1210), .A2(new_n457), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(G50), .C2(new_n801), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n782), .A2(new_n771), .B1(new_n790), .B2(new_n342), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n789), .A2(new_n1175), .B1(new_n770), .B2(new_n1197), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n776), .A2(new_n622), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n782), .A2(new_n218), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n789), .A2(new_n525), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n770), .A2(new_n848), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n787), .A2(new_n805), .B1(new_n790), .B2(new_n498), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1267), .A2(new_n1031), .A3(new_n1066), .A4(new_n457), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1258), .A2(new_n1261), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1255), .B1(new_n844), .B2(new_n1269), .C1(new_n929), .C2(new_n762), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(KEYINPUT121), .B1(new_n1254), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT121), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n1270), .C1(new_n1161), .C2(new_n747), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1253), .A2(new_n1275), .ZN(G381));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1279), .A2(G387), .A3(G381), .A4(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G407));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT122), .Z(new_n1286));
  OAI21_X1  g1086(.A(new_n1282), .B1(new_n1281), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(G213), .ZN(G409));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(G378), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1285), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1119), .A2(new_n1130), .A3(new_n1151), .A4(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n690), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT60), .B1(new_n1161), .B2(new_n1151), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1252), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1278), .B1(new_n1292), .B2(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1293), .A2(new_n690), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1252), .B1(new_n1163), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1275), .A3(G384), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1251), .B(new_n1244), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1243), .A2(new_n1169), .A3(new_n1193), .A4(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1290), .A2(new_n1291), .A3(new_n1304), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n748), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1305), .A2(new_n1310), .A3(new_n1226), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(G378), .A2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(G378), .B2(G375), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1286), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1314), .A4(new_n1304), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1309), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT125), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1290), .A2(new_n1314), .A3(new_n1306), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1286), .A2(G2897), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1301), .A2(new_n1275), .A3(G384), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1301), .B2(new_n1275), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1319), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1285), .A2(G2897), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1297), .A2(new_n1302), .A3(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1322), .A2(new_n1324), .A3(KEYINPUT123), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT123), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1303), .A2(new_n1326), .A3(new_n1319), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1318), .B2(new_n1328), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1316), .A2(new_n1317), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1317), .B1(new_n1316), .B2(new_n1329), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(G393), .B(new_n815), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1017), .A2(new_n1041), .A3(G390), .ZN(new_n1334));
  AOI21_X1  g1134(.A(G390), .B1(new_n1017), .B2(new_n1041), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1333), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G387), .A2(new_n1277), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1017), .A2(new_n1041), .A3(G390), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1332), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1340), .A2(KEYINPUT126), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(KEYINPUT126), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1330), .A2(new_n1331), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1310), .A2(new_n1226), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1151), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1347), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n691), .B1(new_n1348), .B2(KEYINPUT57), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1244), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT57), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1346), .B1(new_n1349), .B2(new_n1352), .ZN(new_n1353));
  AOI211_X1 g1153(.A(KEYINPUT117), .B(new_n691), .C1(new_n1156), .C2(new_n1163), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1167), .B1(new_n1153), .B2(new_n690), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1192), .B1(new_n1356), .B2(new_n1166), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1291), .B(new_n1306), .C1(new_n1353), .C2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1328), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(KEYINPUT63), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1307), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT61), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1336), .A2(new_n1339), .A3(new_n1362), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1290), .A2(new_n1314), .A3(new_n1304), .A4(new_n1306), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1363), .B1(new_n1365), .B2(KEYINPUT63), .ZN(new_n1366));
  AOI21_X1  g1166(.A(KEYINPUT124), .B1(new_n1361), .B2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1352), .A2(new_n690), .A3(new_n1247), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1357), .B1(new_n1368), .B2(new_n1243), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1369), .A2(new_n1285), .A3(new_n1312), .ZN(new_n1370));
  AOI22_X1  g1170(.A1(new_n1359), .A2(KEYINPUT63), .B1(new_n1370), .B2(new_n1304), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT124), .ZN(new_n1372));
  AND3_X1   g1172(.A1(new_n1336), .A2(new_n1339), .A3(new_n1362), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1373), .B1(new_n1364), .B2(new_n1374), .ZN(new_n1375));
  NOR3_X1   g1175(.A1(new_n1371), .A2(new_n1372), .A3(new_n1375), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1367), .A2(new_n1376), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1289), .B1(new_n1345), .B2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1361), .A2(KEYINPUT124), .A3(new_n1366), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1372), .B1(new_n1371), .B2(new_n1375), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  AND2_X1   g1181(.A1(new_n1316), .A2(new_n1329), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1343), .B1(new_n1382), .B2(new_n1317), .ZN(new_n1383));
  OAI211_X1 g1183(.A(KEYINPUT127), .B(new_n1381), .C1(new_n1383), .C2(new_n1330), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1378), .A2(new_n1384), .ZN(G405));
  NOR2_X1   g1185(.A1(new_n1282), .A2(new_n1369), .ZN(new_n1386));
  XNOR2_X1  g1186(.A(new_n1386), .B(new_n1304), .ZN(new_n1387));
  XNOR2_X1  g1187(.A(new_n1387), .B(new_n1340), .ZN(G402));
endmodule


