//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1243,
    new_n1244, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT65), .Z(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G107), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G50), .B2(G226), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n209), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  AND2_X1   g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n204), .A2(G50), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n221), .B(new_n224), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G20), .ZN(new_n249));
  AND3_X1   g0049(.A1(new_n249), .A2(KEYINPUT69), .A3(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(KEYINPUT69), .B1(new_n249), .B2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(new_n210), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n255), .A2(new_n256), .B1(new_n249), .B2(G68), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n248), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT11), .ZN(new_n259));
  INV_X1    g0059(.A(new_n248), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT68), .B(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(new_n249), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT12), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n261), .A2(new_n264), .A3(new_n249), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n265), .B2(new_n203), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G13), .A3(G20), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n259), .B1(new_n203), .B2(new_n262), .C1(new_n266), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G226), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(G232), .A3(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G97), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n279), .B(new_n280), .C1(new_n254), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G41), .A2(G45), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n284), .B1(new_n261), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n282), .A2(new_n285), .B1(G238), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n286), .A2(G1), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n289), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n276), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(G169), .A3(new_n275), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n294), .A2(G179), .A3(new_n296), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n303), .B(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n274), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n274), .B1(new_n297), .B2(G200), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n298), .A2(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n310));
  INV_X1    g0110(.A(G150), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT8), .B(G58), .Z(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n310), .B1(new_n311), .B2(new_n255), .C1(new_n313), .C2(new_n252), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(new_n248), .B1(new_n256), .B2(new_n265), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n262), .A2(new_n256), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G226), .ZN(new_n318));
  MUX2_X1   g0118(.A(G222), .B(G223), .S(G1698), .Z(new_n319));
  NAND2_X1  g0119(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G33), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n285), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n277), .A2(G77), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n292), .B1(new_n287), .B2(new_n318), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n299), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n317), .B(new_n327), .C1(G179), .C2(new_n326), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n277), .A2(G238), .A3(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n212), .C2(new_n277), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n331), .A2(KEYINPUT70), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(KEYINPUT70), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n285), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n291), .B1(new_n288), .B2(G244), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G13), .A2(G33), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(new_n207), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n210), .B1(new_n262), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n255), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n312), .A3(new_n343), .ZN(new_n344));
  XOR2_X1   g0144(.A(KEYINPUT15), .B(G87), .Z(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n251), .B2(new_n250), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n248), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G77), .B2(new_n272), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(G169), .B1(new_n334), .B2(new_n335), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n337), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n306), .A2(new_n309), .A3(new_n328), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n326), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n326), .A2(G200), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  AND3_X1   g0159(.A1(new_n315), .A2(new_n359), .A3(new_n316), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n315), .B2(new_n316), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n357), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(KEYINPUT72), .A2(KEYINPUT10), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n355), .A3(new_n363), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n349), .B1(new_n336), .B2(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n356), .B2(new_n336), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G232), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n292), .B1(new_n287), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n320), .A2(new_n322), .A3(G223), .A4(new_n278), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT77), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n277), .A2(KEYINPUT77), .A3(G223), .A4(new_n278), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n277), .A2(G226), .A3(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n371), .B1(new_n378), .B2(new_n285), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n379), .A2(G179), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n299), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT78), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n204), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n341), .A2(G159), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(KEYINPUT75), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n249), .B1(new_n204), .B2(new_n384), .ZN(new_n390));
  INV_X1    g0190(.A(G159), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n255), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n254), .A3(KEYINPUT3), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(G20), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n398), .C1(new_n323), .C2(new_n395), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n277), .B2(G20), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n203), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n383), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n323), .A2(new_n398), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n323), .B2(new_n249), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n393), .A4(new_n388), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(new_n406), .A3(new_n248), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n262), .A2(new_n312), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n265), .B2(new_n312), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n379), .A2(G179), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n412), .C1(new_n299), .C2(new_n379), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n382), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n379), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n379), .A2(G190), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n418), .A2(new_n407), .A3(new_n409), .A4(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  NOR2_X1   g0223(.A1(KEYINPUT79), .A2(KEYINPUT18), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n415), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n382), .A2(new_n410), .A3(new_n413), .A4(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n416), .A2(new_n422), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n354), .A2(new_n369), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n290), .B1(new_n225), .B2(new_n283), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT5), .B(G41), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n271), .A2(new_n430), .A3(G45), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n213), .A2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G257), .B2(G1698), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n284), .B1(new_n433), .B2(new_n277), .ZN(new_n434));
  INV_X1    g0234(.A(G303), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n323), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n429), .A2(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G45), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n268), .B2(new_n270), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n430), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(G270), .A3(new_n284), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n299), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n265), .A2(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n246), .A2(new_n247), .B1(G20), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G283), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n249), .C1(G33), .C2(new_n281), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n445), .A2(KEYINPUT20), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT20), .B1(new_n445), .B2(new_n447), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n271), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n272), .A2(new_n260), .A3(new_n450), .ZN(new_n451));
  OAI221_X1 g0251(.A(new_n444), .B1(new_n448), .B2(new_n449), .C1(new_n451), .C2(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT21), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n434), .A2(new_n436), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n439), .A2(new_n429), .A3(new_n430), .ZN(new_n456));
  AND4_X1   g0256(.A1(G179), .A2(new_n441), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n453), .A2(new_n454), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT86), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n453), .B2(new_n454), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n442), .A2(KEYINPUT86), .A3(new_n452), .A4(KEYINPUT21), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n272), .A2(new_n345), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT19), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT83), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT83), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT19), .ZN(new_n467));
  AND2_X1   g0267(.A1(G33), .A2(G97), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n249), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(G87), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G97), .B1(new_n250), .B2(new_n251), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n465), .A2(new_n467), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n277), .A2(new_n249), .A3(G68), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n463), .B1(new_n481), .B2(new_n248), .ZN(new_n482));
  INV_X1    g0282(.A(new_n451), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n345), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n429), .A2(new_n261), .A3(new_n438), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n271), .A2(G45), .B1(new_n284), .B2(G250), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT82), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(G33), .A2(G41), .ZN(new_n489));
  OAI21_X1  g0289(.A(G250), .B1(new_n489), .B2(new_n247), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n261), .B2(new_n438), .ZN(new_n491));
  OAI21_X1  g0291(.A(G274), .B1(new_n489), .B2(new_n247), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n439), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n211), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n277), .B(new_n496), .C1(G238), .C2(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n488), .A2(new_n495), .B1(new_n285), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G179), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n485), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n500), .A2(G169), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n285), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n494), .B1(new_n491), .B2(new_n493), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(G190), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT85), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n451), .B2(new_n472), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n249), .B1(new_n268), .B2(new_n270), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n248), .B1(new_n511), .B2(G13), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(KEYINPUT85), .A3(G87), .A4(new_n450), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n482), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n500), .A2(new_n417), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n503), .A2(new_n504), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n452), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n441), .A2(new_n455), .A3(new_n456), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n437), .A2(G190), .A3(new_n441), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n417), .B1(new_n437), .B2(new_n441), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT87), .B1(new_n524), .B2(new_n452), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n462), .A2(new_n517), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n212), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n272), .B2(G107), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n483), .A2(G107), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n320), .A2(new_n322), .A3(new_n249), .A4(G87), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(KEYINPUT88), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n277), .A2(new_n249), .A3(G87), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT23), .B1(new_n249), .B2(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT89), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT89), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(KEYINPUT23), .C1(new_n249), .C2(G107), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n498), .A2(G20), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n249), .A2(KEYINPUT23), .A3(G107), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT24), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n545), .B(new_n543), .C1(new_n539), .C2(new_n541), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n534), .A4(new_n536), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT90), .B1(new_n552), .B2(new_n248), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT90), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n554), .B(new_n260), .C1(new_n548), .C2(new_n551), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n531), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g0356(.A1(G250), .A2(G1698), .ZN(new_n557));
  INV_X1    g0357(.A(G257), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G1698), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n320), .A2(new_n557), .A3(new_n322), .A4(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(new_n254), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n285), .B1(new_n439), .B2(new_n430), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n285), .A2(new_n562), .B1(new_n563), .B2(G264), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n564), .A2(new_n456), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G179), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n285), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT91), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n563), .A2(G264), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(KEYINPUT91), .A3(new_n285), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n569), .A2(new_n456), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G169), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n556), .A2(new_n574), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n565), .A2(G200), .B1(new_n572), .B2(G190), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(new_n531), .C1(new_n553), .C2(new_n555), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(G257), .A2(new_n563), .B1(new_n431), .B2(new_n429), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n211), .A2(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(new_n320), .A3(new_n322), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n320), .A2(new_n322), .A3(G250), .A4(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n581), .A2(new_n320), .A3(new_n322), .A4(KEYINPUT4), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n584), .A2(new_n446), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n285), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n580), .A2(new_n588), .A3(KEYINPUT80), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT80), .B1(new_n580), .B2(new_n588), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(G169), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n399), .A2(new_n400), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n212), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n281), .A2(new_n212), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(new_n471), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(KEYINPUT6), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n592), .A2(G107), .B1(G20), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n341), .A2(G77), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n260), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n265), .A2(new_n281), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n451), .B2(new_n281), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n580), .A2(new_n588), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n599), .A2(new_n601), .B1(G179), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT81), .B1(new_n591), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n592), .A2(G107), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n596), .A2(G20), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n598), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n601), .B1(new_n607), .B2(new_n248), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n602), .A2(G179), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n580), .A2(new_n588), .A3(KEYINPUT80), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n299), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n613), .A2(new_n614), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(G190), .B1(G200), .B2(new_n602), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n604), .A2(new_n616), .B1(new_n608), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n428), .A2(new_n527), .A3(new_n579), .A4(new_n619), .ZN(G372));
  INV_X1    g0420(.A(KEYINPUT94), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n423), .A2(new_n422), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n309), .A2(new_n352), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n306), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n411), .B1(new_n299), .B2(new_n379), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n410), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT18), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n621), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT95), .ZN(new_n629));
  INV_X1    g0429(.A(new_n366), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(new_n364), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n365), .A2(KEYINPUT95), .A3(new_n366), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT18), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n626), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n303), .B(KEYINPUT74), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n300), .A3(new_n301), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n274), .B1(new_n309), .B2(new_n352), .ZN(new_n638));
  OAI211_X1 g0438(.A(KEYINPUT94), .B(new_n635), .C1(new_n638), .C2(new_n622), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n328), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n642));
  INV_X1    g0442(.A(new_n556), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(new_n575), .B1(new_n643), .B2(new_n576), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT92), .B1(new_n506), .B2(new_n507), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT92), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n488), .A2(new_n495), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n505), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n299), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n482), .A2(new_n484), .B1(new_n500), .B2(new_n501), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n515), .B1(G200), .B2(new_n648), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT93), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n650), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n648), .A2(G200), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n508), .A2(new_n482), .A3(new_n514), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n644), .A2(new_n660), .A3(new_n619), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n591), .A2(new_n603), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n654), .B2(new_n657), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n504), .ZN(new_n667));
  INV_X1    g0467(.A(new_n516), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n667), .A2(new_n650), .B1(new_n668), .B2(new_n656), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n604), .A3(new_n616), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT26), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n661), .A2(new_n654), .A3(new_n666), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n428), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n641), .A2(new_n673), .ZN(G369));
  NOR2_X1   g0474(.A1(new_n264), .A2(G20), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n261), .A2(new_n676), .A3(KEYINPUT27), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT27), .B1(new_n261), .B2(new_n676), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(G213), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n643), .A2(new_n682), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n578), .A2(new_n683), .B1(new_n575), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n462), .A2(new_n682), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n518), .A2(new_n682), .ZN(new_n689));
  OR3_X1    g0489(.A1(new_n462), .A2(new_n526), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n462), .A2(new_n689), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n556), .A2(new_n574), .A3(new_n682), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n579), .A2(new_n686), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n222), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G1), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n473), .A2(new_n474), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n443), .A3(new_n471), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n700), .A2(new_n702), .B1(new_n227), .B2(new_n699), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT98), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT97), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n589), .A2(new_n590), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n500), .A2(new_n457), .A3(new_n564), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n709), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n456), .A2(new_n564), .B1(new_n580), .B2(new_n588), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n648), .A2(new_n714), .A3(new_n501), .A4(new_n520), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n564), .A2(G179), .A3(new_n437), .A4(new_n441), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n505), .B(new_n711), .C1(new_n506), .C2(new_n507), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n617), .A2(new_n718), .A3(new_n708), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n713), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n721));
  AND3_X1   g0521(.A1(new_n720), .A2(new_n681), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n720), .B2(new_n681), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n705), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n720), .A2(new_n681), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n720), .A2(new_n681), .A3(new_n721), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(KEYINPUT98), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n579), .A2(new_n619), .A3(new_n527), .A4(new_n682), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT99), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n731), .A2(new_n732), .A3(G330), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(new_n731), .B2(G330), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT26), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n670), .A2(new_n662), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(KEYINPUT100), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT100), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n660), .A2(new_n740), .A3(KEYINPUT26), .A4(new_n663), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n739), .A2(new_n654), .A3(new_n661), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n736), .B1(new_n742), .B2(new_n682), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n672), .A2(new_n736), .A3(new_n682), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n735), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n704), .B1(new_n747), .B2(G1), .ZN(G364));
  XOR2_X1   g0548(.A(new_n692), .B(KEYINPUT101), .Z(new_n749));
  AOI21_X1  g0549(.A(new_n267), .B1(new_n675), .B2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n698), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n690), .A2(new_n691), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n749), .B(new_n753), .C1(G330), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n249), .A2(new_n501), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G200), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G311), .A2(new_n758), .B1(new_n760), .B2(G322), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G20), .A3(new_n356), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G329), .ZN(new_n765));
  INV_X1    g0565(.A(G326), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n759), .A2(new_n417), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n761), .B(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n757), .A2(new_n417), .A3(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OR2_X1    g0571(.A1(KEYINPUT33), .A2(G317), .ZN(new_n772));
  NAND2_X1  g0572(.A1(KEYINPUT33), .A2(G317), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n249), .A2(new_n417), .A3(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n356), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n769), .A2(new_n277), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n762), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n775), .A2(G190), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT105), .ZN(new_n784));
  OAI221_X1 g0584(.A(new_n779), .B1(new_n561), .B2(new_n782), .C1(new_n435), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT106), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n771), .A2(new_n203), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(new_n281), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n277), .B1(new_n768), .B2(new_n256), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT32), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT104), .B(G159), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n764), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n776), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G107), .ZN(new_n796));
  INV_X1    g0596(.A(new_n760), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n797), .B2(new_n202), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n793), .A2(new_n790), .B1(new_n701), .B2(new_n783), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n758), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n794), .B(new_n800), .C1(new_n210), .C2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n786), .B1(new_n787), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n247), .B1(G20), .B2(new_n299), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n338), .B(KEYINPUT102), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n249), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT103), .Z(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n804), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n277), .A2(G355), .A3(new_n222), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n697), .A2(new_n277), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n244), .B2(new_n438), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n227), .A2(G45), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n810), .B1(G116), .B2(new_n222), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n803), .A2(new_n804), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n815), .B(new_n752), .C1(new_n754), .C2(new_n807), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n755), .A2(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n352), .A2(new_n682), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n368), .B1(new_n350), .B2(new_n682), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n353), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n735), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n733), .B2(new_n734), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n672), .A2(new_n682), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n825), .B(new_n826), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n753), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n758), .A2(new_n791), .B1(new_n760), .B2(G143), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n829), .B1(new_n830), .B2(new_n768), .C1(new_n311), .C2(new_n771), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(new_n784), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(G50), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n781), .A2(G58), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n323), .B1(new_n764), .B2(G132), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n795), .A2(G68), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n843), .A2(new_n777), .B1(new_n443), .B2(new_n801), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT108), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(new_n435), .C2(new_n768), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT109), .Z(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n323), .B1(new_n763), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n851), .B(new_n788), .C1(G294), .C2(new_n760), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n849), .B(new_n852), .C1(new_n472), .C2(new_n776), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n784), .A2(new_n212), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n804), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n822), .A2(new_n805), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n804), .A2(new_n338), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n210), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n856), .A2(new_n752), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n828), .A2(new_n860), .ZN(G384));
  NAND3_X1  g0661(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n726), .A2(new_n721), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n730), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n821), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n274), .A2(new_n681), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n306), .A2(new_n309), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n637), .A2(new_n274), .A3(new_n681), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT110), .ZN(new_n871));
  INV_X1    g0671(.A(new_n679), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n410), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n626), .A2(new_n873), .A3(new_n420), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n874), .B2(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n414), .A2(new_n877), .A3(new_n420), .A4(new_n873), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n874), .A2(new_n871), .A3(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n420), .B(KEYINPUT17), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n873), .B1(new_n635), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n406), .A2(new_n248), .ZN(new_n885));
  INV_X1    g0685(.A(new_n394), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n886), .B2(new_n405), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n409), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n872), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n427), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n625), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n889), .A2(new_n892), .A3(new_n420), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT40), .B1(new_n870), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n891), .B2(new_n895), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n865), .A4(new_n869), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n428), .A2(new_n864), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT39), .B1(new_n896), .B2(new_n899), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n874), .A2(new_n871), .A3(KEYINPUT37), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n875), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n882), .B1(new_n913), .B2(new_n878), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n915), .B2(KEYINPUT39), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n637), .A2(new_n274), .A3(new_n682), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n867), .A2(new_n868), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n820), .A2(new_n353), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n672), .A2(new_n682), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n922), .B2(new_n818), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n900), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n627), .A2(new_n679), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n909), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n428), .B1(new_n743), .B2(new_n744), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n641), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n271), .B2(new_n675), .ZN(new_n932));
  OAI211_X1 g0732(.A(G20), .B(new_n225), .C1(new_n596), .C2(KEYINPUT35), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n443), .B(new_n933), .C1(KEYINPUT35), .C2(new_n596), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT36), .Z(new_n935));
  AOI211_X1 g0735(.A(new_n210), .B(new_n227), .C1(G58), .C2(G68), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n201), .A2(new_n203), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n264), .B(new_n261), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n932), .A2(new_n935), .A3(new_n938), .ZN(G367));
  OAI22_X1  g0739(.A1(new_n801), .A2(new_n777), .B1(new_n797), .B2(new_n435), .ZN(new_n940));
  INV_X1    g0740(.A(new_n843), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(G294), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT46), .B1(new_n784), .B2(new_n443), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n783), .A2(KEYINPUT46), .A3(new_n443), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n767), .A2(G311), .B1(G107), .B2(new_n781), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n776), .A2(new_n281), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n277), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n940), .B(new_n949), .C1(G317), .C2(new_n764), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n783), .A2(new_n202), .B1(new_n830), .B2(new_n763), .ZN(new_n951));
  INV_X1    g0751(.A(new_n201), .ZN(new_n952));
  INV_X1    g0752(.A(G143), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n801), .A2(new_n952), .B1(new_n768), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G68), .B2(new_n781), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n323), .B1(new_n795), .B2(G77), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(new_n311), .C2(new_n797), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n951), .B(new_n957), .C1(new_n791), .C2(new_n941), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT114), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT47), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n804), .ZN(new_n962));
  INV_X1    g0762(.A(new_n345), .ZN(new_n963));
  INV_X1    g0763(.A(new_n811), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n809), .B1(new_n222), .B2(new_n963), .C1(new_n237), .C2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n752), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n482), .A2(new_n514), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n681), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n654), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n660), .B2(new_n968), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n970), .A2(new_n808), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT43), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n604), .A2(new_n616), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n619), .B1(new_n608), .B2(new_n682), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n663), .A2(new_n681), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n975), .B1(new_n979), .B2(new_n575), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT111), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n682), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n695), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT42), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n974), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n970), .A2(new_n973), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n693), .A2(new_n979), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n987), .A2(new_n988), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n995), .B2(new_n989), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n695), .A2(new_n694), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n979), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n979), .A2(new_n998), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(new_n693), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT112), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n693), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n687), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n749), .B1(new_n984), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(new_n747), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n747), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n698), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n751), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT113), .B1(new_n997), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n994), .A2(new_n996), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT113), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1014), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n1012), .B2(new_n747), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1017), .B(new_n1018), .C1(new_n751), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n972), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n1011), .A2(new_n747), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n699), .B1(new_n1010), .B2(new_n746), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n782), .A2(new_n777), .B1(new_n783), .B2(new_n561), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT115), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G303), .A2(new_n758), .B1(new_n760), .B2(G317), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n767), .A2(G322), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n843), .C2(new_n850), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1028), .B1(new_n1032), .B2(KEYINPUT48), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(KEYINPUT115), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT116), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT48), .B2(new_n1032), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT49), .Z(new_n1038));
  OAI22_X1  g0838(.A1(new_n776), .A2(new_n443), .B1(new_n766), .B2(new_n763), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n277), .A3(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n801), .A2(new_n203), .B1(new_n210), .B2(new_n783), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n312), .B2(new_n770), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n256), .B2(new_n797), .C1(new_n311), .C2(new_n763), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n277), .B1(new_n782), .B2(new_n963), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n768), .A2(new_n391), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1043), .A2(new_n947), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n804), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n684), .A2(new_n807), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n312), .A2(new_n256), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n203), .A2(new_n210), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1050), .A2(G45), .A3(new_n1051), .A4(new_n702), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n811), .B1(new_n234), .B2(new_n438), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n702), .A2(new_n222), .A3(new_n277), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n222), .A2(G107), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n809), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1047), .A2(new_n752), .A3(new_n1048), .A4(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1026), .B(new_n1058), .C1(new_n750), .C2(new_n1010), .ZN(G393));
  INV_X1    g0859(.A(new_n693), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1004), .B(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(KEYINPUT118), .A3(new_n1024), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(new_n1012), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT118), .B1(new_n1061), .B2(new_n1024), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1064), .A2(new_n699), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT119), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT119), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1005), .A2(new_n751), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n753), .B1(new_n979), .B2(new_n808), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n809), .B1(new_n281), .B2(new_n222), .C1(new_n241), .C2(new_n964), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G150), .A2(new_n767), .B1(new_n760), .B2(G159), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n472), .B2(new_n776), .C1(new_n952), .C2(new_n843), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n763), .A2(new_n953), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n801), .A2(new_n313), .B1(new_n210), .B2(new_n782), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n277), .B1(new_n783), .B2(new_n203), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n796), .B1(new_n777), .B2(new_n783), .C1(new_n843), .C2(new_n435), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n767), .A2(G317), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n797), .B2(new_n850), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n277), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n758), .A2(G294), .B1(G116), .B2(new_n781), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1081), .B(new_n1087), .C1(G322), .C2(new_n764), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n804), .B1(new_n1080), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1072), .A2(new_n1073), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1070), .A2(new_n1071), .A3(new_n1090), .ZN(G390));
  OAI211_X1 g0891(.A(new_n821), .B(new_n869), .C1(new_n733), .C2(new_n734), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n865), .A2(G330), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n920), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n742), .A2(new_n682), .A3(new_n921), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n818), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n865), .A2(G330), .A3(new_n869), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n824), .B2(new_n920), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n922), .A2(new_n818), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n641), .A2(new_n906), .A3(new_n929), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1101), .A2(new_n869), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n916), .B1(new_n1107), .B2(new_n917), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n915), .A2(new_n917), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1096), .B2(new_n869), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1108), .A2(new_n1110), .B1(new_n688), .B2(new_n870), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1096), .A2(new_n869), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1109), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1092), .ZN(new_n1115));
  OR3_X1    g0915(.A1(new_n884), .A2(new_n896), .A3(KEYINPUT39), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n910), .B(new_n1116), .C1(new_n923), .C2(new_n918), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1106), .A2(new_n1111), .A3(new_n1118), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1108), .A2(new_n1092), .A3(new_n1110), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1099), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1103), .B(new_n1105), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n750), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1116), .A2(new_n805), .A3(new_n910), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G294), .A2(new_n764), .B1(new_n781), .B2(G77), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n323), .C1(new_n768), .C2(new_n777), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n835), .A2(G87), .B1(G116), .B2(new_n760), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1128), .B(new_n839), .C1(new_n212), .C2(new_n843), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(G97), .C2(new_n758), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n941), .A2(G137), .B1(G132), .B2(new_n760), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n768), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT53), .B1(new_n783), .B2(new_n311), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1134), .B(new_n277), .C1(new_n391), .C2(new_n782), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n311), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n795), .A2(new_n201), .B1(G125), .B2(new_n764), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1137), .B1(new_n801), .B2(new_n1139), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .A4(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n804), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n858), .A2(new_n313), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1125), .A2(new_n752), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OR3_X1    g0945(.A1(new_n1124), .A2(KEYINPUT120), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT120), .B1(new_n1124), .B2(new_n1145), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1123), .A2(new_n698), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  NAND2_X1  g0949(.A1(new_n317), .A2(new_n872), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n631), .A2(new_n632), .A3(new_n328), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(KEYINPUT122), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT122), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n631), .A2(new_n632), .A3(new_n1153), .A4(new_n328), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1150), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n1154), .A3(new_n1150), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1157), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1152), .A2(new_n1154), .A3(new_n1150), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n1155), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(new_n903), .A3(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n903), .B2(G330), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n926), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n904), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n927), .A3(new_n1164), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n751), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1163), .A2(new_n805), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n770), .A2(G132), .B1(new_n767), .B2(G125), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n758), .A2(G137), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n783), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1175), .A2(new_n1138), .B1(new_n781), .B2(G150), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G128), .B2(new_n760), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G33), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n795), .A2(new_n791), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G41), .B1(new_n764), .B2(G124), .ZN(new_n1183));
  AND4_X1   g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n797), .A2(new_n212), .B1(new_n203), .B2(new_n782), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n776), .A2(new_n202), .B1(new_n777), .B2(new_n763), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n783), .A2(new_n210), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1186), .A2(new_n1187), .A3(G41), .A4(new_n277), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT121), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1185), .B(new_n1189), .C1(new_n345), .C2(new_n758), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n281), .B2(new_n771), .C1(new_n443), .C2(new_n768), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .C1(G50), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n804), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n858), .A2(new_n952), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1172), .A2(new_n752), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1171), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1104), .B(KEYINPUT123), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1122), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT124), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1122), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1201), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n698), .B1(new_n1207), .B2(KEYINPUT57), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1122), .A2(KEYINPUT124), .A3(new_n1202), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT124), .B1(new_n1122), .B2(new_n1202), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1170), .B(KEYINPUT57), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1200), .B1(new_n1208), .B2(new_n1212), .ZN(G375));
  OR2_X1    g1013(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1014), .A3(new_n1106), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n920), .A2(new_n338), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n277), .B1(new_n763), .B2(new_n1132), .C1(new_n801), .C2(new_n311), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G132), .A2(new_n767), .B1(new_n760), .B2(G137), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n843), .B2(new_n1139), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT125), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n256), .B2(new_n782), .C1(new_n202), .C2(new_n776), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1217), .B(new_n1221), .C1(G159), .C2(new_n835), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n835), .A2(G97), .B1(G294), .B2(new_n767), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n443), .B2(new_n843), .C1(new_n777), .C2(new_n797), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n763), .A2(new_n435), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n323), .B1(new_n776), .B2(new_n210), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n801), .A2(new_n212), .B1(new_n963), .B2(new_n782), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n804), .B1(new_n1222), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n858), .A2(new_n203), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1216), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1103), .A2(new_n751), .B1(new_n752), .B2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1215), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G381));
  NAND4_X1  g1034(.A1(new_n1022), .A2(new_n1071), .A3(new_n1070), .A4(new_n1090), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G396), .A3(G393), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1123), .A2(new_n698), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1124), .A2(new_n1145), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(G375), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1236), .A2(new_n1237), .A3(new_n1233), .A4(new_n1241), .ZN(G407));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1241), .B2(new_n680), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G407), .A2(new_n1244), .ZN(G409));
  OAI21_X1  g1045(.A(new_n1170), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT57), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n699), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1148), .B(new_n1199), .C1(new_n1248), .C2(new_n1211), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1207), .A2(new_n1014), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1240), .B1(new_n1200), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT126), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1214), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1214), .A2(new_n1253), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n698), .A3(new_n1106), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1232), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1237), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(G384), .A3(new_n1232), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1243), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1251), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1200), .C1(new_n1208), .C2(new_n1212), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1252), .A2(new_n1260), .A3(new_n1262), .A4(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1259), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1261), .B(new_n1270), .C1(new_n1264), .C2(new_n1263), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT61), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1261), .A2(G2897), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1260), .B(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1261), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1275), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1273), .A2(new_n1274), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(G390), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1235), .ZN(new_n1283));
  XOR2_X1   g1083(.A(G393), .B(G396), .Z(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1282), .A2(new_n1235), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1271), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1279), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1281), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1278), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1288), .B1(new_n1260), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1267), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1277), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1252), .A2(new_n1262), .A3(new_n1266), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1293), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1295), .B(new_n1275), .C1(new_n1296), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1291), .A2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(new_n1240), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1249), .B1(G375), .B2(new_n1302), .ZN(new_n1303));
  XOR2_X1   g1103(.A(new_n1303), .B(new_n1260), .Z(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1288), .ZN(G402));
endmodule


