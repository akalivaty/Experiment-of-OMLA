

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575;

  XNOR2_X1 U321 ( .A(n340), .B(KEYINPUT33), .ZN(n341) );
  XNOR2_X1 U322 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U323 ( .A(n404), .B(KEYINPUT48), .ZN(n536) );
  XNOR2_X1 U324 ( .A(n446), .B(G176GAT), .ZN(n447) );
  XNOR2_X1 U325 ( .A(n448), .B(n447), .ZN(G1349GAT) );
  XOR2_X1 U326 ( .A(KEYINPUT17), .B(KEYINPUT79), .Z(n290) );
  XNOR2_X1 U327 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n289) );
  XNOR2_X1 U328 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U329 ( .A(KEYINPUT19), .B(n291), .Z(n418) );
  XOR2_X1 U330 ( .A(KEYINPUT20), .B(KEYINPUT78), .Z(n293) );
  XNOR2_X1 U331 ( .A(G169GAT), .B(KEYINPUT81), .ZN(n292) );
  XNOR2_X1 U332 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U333 ( .A(G71GAT), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U334 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U336 ( .A(n297), .B(n296), .Z(n308) );
  XOR2_X1 U337 ( .A(G127GAT), .B(G134GAT), .Z(n299) );
  XNOR2_X1 U338 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U339 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U340 ( .A(G113GAT), .B(n300), .Z(n442) );
  XOR2_X1 U341 ( .A(KEYINPUT82), .B(G190GAT), .Z(n302) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .ZN(n301) );
  XNOR2_X1 U343 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U344 ( .A(KEYINPUT77), .B(n303), .Z(n305) );
  NAND2_X1 U345 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U346 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n442), .B(n306), .ZN(n307) );
  XNOR2_X1 U348 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U349 ( .A(n418), .B(n309), .Z(n460) );
  INV_X1 U350 ( .A(n460), .ZN(n518) );
  NAND2_X1 U351 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U352 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n311) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(KEYINPUT88), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U355 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n312) );
  XNOR2_X1 U356 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U357 ( .A(n315), .B(n314), .ZN(n324) );
  XOR2_X1 U358 ( .A(KEYINPUT87), .B(KEYINPUT83), .Z(n322) );
  XOR2_X1 U359 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U360 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n316) );
  XNOR2_X1 U361 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U362 ( .A(G197GAT), .B(n318), .Z(n409) );
  XOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT69), .Z(n320) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n320), .B(n319), .ZN(n375) );
  XNOR2_X1 U366 ( .A(n409), .B(n375), .ZN(n321) );
  XNOR2_X1 U367 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U368 ( .A(n324), .B(n323), .ZN(n330) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT2), .Z(n326) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n325) );
  XNOR2_X1 U371 ( .A(n326), .B(n325), .ZN(n436) );
  XOR2_X1 U372 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U373 ( .A(G106GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n337) );
  XNOR2_X1 U375 ( .A(n436), .B(n337), .ZN(n329) );
  XNOR2_X1 U376 ( .A(n330), .B(n329), .ZN(n459) );
  XOR2_X1 U377 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n423) );
  XOR2_X1 U378 ( .A(G71GAT), .B(G57GAT), .Z(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT13), .B(n331), .Z(n360) );
  XOR2_X1 U380 ( .A(KEYINPUT67), .B(KEYINPUT32), .Z(n333) );
  NAND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(n334), .B(KEYINPUT31), .Z(n339) );
  XOR2_X1 U384 ( .A(KEYINPUT68), .B(G92GAT), .Z(n336) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n374) );
  XNOR2_X1 U387 ( .A(n337), .B(n374), .ZN(n338) );
  XOR2_X1 U388 ( .A(n339), .B(n338), .Z(n342) );
  XOR2_X1 U389 ( .A(G176GAT), .B(G64GAT), .Z(n407) );
  XNOR2_X1 U390 ( .A(G120GAT), .B(n407), .ZN(n340) );
  XOR2_X1 U391 ( .A(n360), .B(n343), .Z(n565) );
  XNOR2_X1 U392 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n379) );
  XOR2_X1 U393 ( .A(G78GAT), .B(G155GAT), .Z(n345) );
  XNOR2_X1 U394 ( .A(G183GAT), .B(G127GAT), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(G64GAT), .Z(n347) );
  XNOR2_X1 U397 ( .A(G8GAT), .B(G211GAT), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U399 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U400 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n351) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U403 ( .A(KEYINPUT12), .B(n352), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U405 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n356) );
  XNOR2_X1 U406 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n358), .B(n357), .Z(n362) );
  XNOR2_X1 U409 ( .A(G15GAT), .B(G22GAT), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n359), .B(G1GAT), .ZN(n386) );
  XNOR2_X1 U411 ( .A(n386), .B(n360), .ZN(n361) );
  XOR2_X1 U412 ( .A(n362), .B(n361), .Z(n528) );
  INV_X1 U413 ( .A(n528), .ZN(n569) );
  XOR2_X1 U414 ( .A(G29GAT), .B(G43GAT), .Z(n364) );
  XNOR2_X1 U415 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n387) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(n387), .Z(n366) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U420 ( .A(n367), .B(KEYINPUT9), .Z(n369) );
  XOR2_X1 U421 ( .A(G36GAT), .B(G190GAT), .Z(n417) );
  XNOR2_X1 U422 ( .A(G106GAT), .B(n417), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT64), .B(KEYINPUT70), .Z(n371) );
  XNOR2_X1 U425 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U427 ( .A(n373), .B(n372), .Z(n377) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U429 ( .A(n377), .B(n376), .Z(n553) );
  XNOR2_X1 U430 ( .A(KEYINPUT36), .B(n553), .ZN(n571) );
  NAND2_X1 U431 ( .A1(n569), .A2(n571), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U433 ( .A1(n565), .A2(n380), .ZN(n395) );
  XOR2_X1 U434 ( .A(KEYINPUT65), .B(G197GAT), .Z(n382) );
  XNOR2_X1 U435 ( .A(G113GAT), .B(G141GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n394) );
  XOR2_X1 U437 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n384) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n385), .B(KEYINPUT29), .Z(n389) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U443 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XOR2_X1 U444 ( .A(n390), .B(n410), .Z(n392) );
  XNOR2_X1 U445 ( .A(G50GAT), .B(G36GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n560) );
  INV_X1 U448 ( .A(n560), .ZN(n520) );
  NAND2_X1 U449 ( .A1(n395), .A2(n520), .ZN(n403) );
  XOR2_X1 U450 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n397) );
  XNOR2_X1 U451 ( .A(KEYINPUT41), .B(n565), .ZN(n523) );
  INV_X1 U452 ( .A(n523), .ZN(n542) );
  NAND2_X1 U453 ( .A1(n542), .A2(n560), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  NOR2_X1 U455 ( .A1(n569), .A2(n398), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(KEYINPUT113), .ZN(n400) );
  NOR2_X1 U457 ( .A1(n553), .A2(n400), .ZN(n401) );
  XNOR2_X1 U458 ( .A(KEYINPUT47), .B(n401), .ZN(n402) );
  NAND2_X1 U459 ( .A1(n403), .A2(n402), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT96), .B(G92GAT), .Z(n406) );
  XNOR2_X1 U461 ( .A(G204GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n414) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U469 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U470 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U471 ( .A(n420), .B(n419), .Z(n507) );
  INV_X1 U472 ( .A(n507), .ZN(n421) );
  NAND2_X1 U473 ( .A1(n536), .A2(n421), .ZN(n422) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n443) );
  XOR2_X1 U475 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n425) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U478 ( .A(KEYINPUT92), .B(n426), .ZN(n440) );
  XOR2_X1 U479 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n428) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(KEYINPUT89), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n430) );
  XNOR2_X1 U483 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n438) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G162GAT), .Z(n434) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G148GAT), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U492 ( .A(n442), .B(n441), .Z(n457) );
  INV_X1 U493 ( .A(n457), .ZN(n505) );
  NAND2_X1 U494 ( .A1(n443), .A2(n505), .ZN(n558) );
  NOR2_X1 U495 ( .A1(n459), .A2(n558), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n444), .B(KEYINPUT55), .ZN(n445) );
  NOR2_X2 U497 ( .A1(n518), .A2(n445), .ZN(n552) );
  NAND2_X1 U498 ( .A1(n552), .A2(n542), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n446) );
  NOR2_X1 U500 ( .A1(n520), .A2(n565), .ZN(n480) );
  NOR2_X1 U501 ( .A1(n518), .A2(n507), .ZN(n449) );
  NOR2_X1 U502 ( .A1(n459), .A2(n449), .ZN(n450) );
  XOR2_X1 U503 ( .A(n450), .B(KEYINPUT98), .Z(n451) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n451), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n453) );
  NAND2_X1 U506 ( .A1(n459), .A2(n518), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n559) );
  XNOR2_X1 U508 ( .A(n507), .B(KEYINPUT27), .ZN(n458) );
  NOR2_X1 U509 ( .A1(n559), .A2(n458), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n455), .A2(n454), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n457), .A2(n456), .ZN(n462) );
  NOR2_X1 U512 ( .A1(n458), .A2(n505), .ZN(n535) );
  XOR2_X1 U513 ( .A(n459), .B(KEYINPUT28), .Z(n513) );
  NAND2_X1 U514 ( .A1(n535), .A2(n513), .ZN(n517) );
  NOR2_X1 U515 ( .A1(n460), .A2(n517), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n477) );
  INV_X1 U517 ( .A(n553), .ZN(n532) );
  NAND2_X1 U518 ( .A1(n569), .A2(n532), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT16), .ZN(n464) );
  XNOR2_X1 U520 ( .A(n464), .B(KEYINPUT76), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n477), .A2(n465), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT99), .B(n466), .Z(n490) );
  NAND2_X1 U523 ( .A1(n480), .A2(n490), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n505), .A2(n474), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT34), .B(n467), .Z(n468) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U527 ( .A1(n507), .A2(n474), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT100), .B(n469), .Z(n470) );
  XNOR2_X1 U529 ( .A(G8GAT), .B(n470), .ZN(G1325GAT) );
  NOR2_X1 U530 ( .A1(n518), .A2(n474), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U533 ( .A(G15GAT), .B(n473), .Z(G1326GAT) );
  NOR2_X1 U534 ( .A1(n513), .A2(n474), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n475), .Z(n476) );
  XNOR2_X1 U536 ( .A(G22GAT), .B(n476), .ZN(G1327GAT) );
  NOR2_X1 U537 ( .A1(n569), .A2(n477), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n571), .A2(n478), .ZN(n479) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(n479), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n504), .A2(n480), .ZN(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT38), .B(n481), .ZN(n488) );
  NOR2_X1 U542 ( .A1(n488), .A2(n505), .ZN(n483) );
  XNOR2_X1 U543 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U545 ( .A(G29GAT), .B(n484), .Z(G1328GAT) );
  NOR2_X1 U546 ( .A1(n488), .A2(n507), .ZN(n485) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n485), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n488), .A2(n518), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT40), .B(n486), .Z(n487) );
  XNOR2_X1 U550 ( .A(G43GAT), .B(n487), .ZN(G1330GAT) );
  NOR2_X1 U551 ( .A1(n513), .A2(n488), .ZN(n489) );
  XOR2_X1 U552 ( .A(G50GAT), .B(n489), .Z(G1331GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n494) );
  NOR2_X1 U554 ( .A1(n560), .A2(n523), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n490), .A2(n503), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n505), .A2(n498), .ZN(n492) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1332GAT) );
  NOR2_X1 U560 ( .A1(n507), .A2(n498), .ZN(n495) );
  XOR2_X1 U561 ( .A(G64GAT), .B(n495), .Z(G1333GAT) );
  NOR2_X1 U562 ( .A1(n518), .A2(n498), .ZN(n496) );
  XOR2_X1 U563 ( .A(KEYINPUT106), .B(n496), .Z(n497) );
  XNOR2_X1 U564 ( .A(G71GAT), .B(n497), .ZN(G1334GAT) );
  NOR2_X1 U565 ( .A1(n498), .A2(n513), .ZN(n502) );
  XOR2_X1 U566 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n500) );
  XNOR2_X1 U567 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n499) );
  XNOR2_X1 U568 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  NAND2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n512) );
  NOR2_X1 U571 ( .A1(n505), .A2(n512), .ZN(n506) );
  XOR2_X1 U572 ( .A(G85GAT), .B(n506), .Z(G1336GAT) );
  NOR2_X1 U573 ( .A1(n507), .A2(n512), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(n510), .ZN(G1337GAT) );
  NOR2_X1 U577 ( .A1(n518), .A2(n512), .ZN(n511) );
  XOR2_X1 U578 ( .A(G99GAT), .B(n511), .Z(G1338GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n515) );
  XNOR2_X1 U580 ( .A(KEYINPUT111), .B(KEYINPUT44), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U584 ( .A1(n536), .A2(n519), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n520), .A2(n531), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1340GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n531), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n527) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n530) );
  NOR2_X1 U594 ( .A1(n528), .A2(n531), .ZN(n529) );
  XOR2_X1 U595 ( .A(n530), .B(n529), .Z(G1342GAT) );
  NOR2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U600 ( .A1(n537), .A2(n559), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT118), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n560), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n541) );
  XNOR2_X1 U605 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n546) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n548), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n569), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n548), .A2(n553), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n560), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U617 ( .A1(n552), .A2(n569), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT58), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G190GAT), .B(n555), .ZN(G1351GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n564) );
  XOR2_X1 U625 ( .A(G197GAT), .B(KEYINPUT59), .Z(n562) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n572) );
  NAND2_X1 U627 ( .A1(n572), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(n564), .B(n563), .Z(G1352GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n567) );
  NAND2_X1 U631 ( .A1(n572), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G204GAT), .B(n568), .ZN(G1353GAT) );
  NAND2_X1 U634 ( .A1(n572), .A2(n569), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n574) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(n575), .ZN(G1355GAT) );
endmodule

