//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  XOR2_X1   g001(.A(G134gat), .B(G162gat), .Z(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT96), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(KEYINPUT89), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT89), .B2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(new_n213), .ZN(new_n215));
  INV_X1    g014(.A(new_n210), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n207), .A2(KEYINPUT15), .B1(new_n216), .B2(new_n209), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n206), .B1(new_n219), .B2(KEYINPUT90), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n221), .B(KEYINPUT17), .C1(new_n214), .C2(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G99gat), .B(G106gat), .Z(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n226), .B(new_n227), .Z(new_n228));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229));
  INV_X1    g028(.A(G85gat), .ZN(new_n230));
  INV_X1    g029(.A(G92gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(KEYINPUT8), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n225), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(new_n225), .A3(new_n232), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT98), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT98), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n238), .ZN(new_n242));
  INV_X1    g041(.A(new_n219), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G232gat), .A2(G233gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT41), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n220), .B2(new_n222), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n246), .ZN(new_n249));
  OAI21_X1  g048(.A(G190gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G218gat), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n205), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n245), .A2(KEYINPUT41), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(G218gat), .A3(new_n250), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n253), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n204), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n254), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n203), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G57gat), .B(G64gat), .Z(new_n265));
  INV_X1    g064(.A(KEYINPUT9), .ZN(new_n266));
  NAND2_X1  g065(.A1(G71gat), .A2(G78gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n265), .A2(KEYINPUT95), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(KEYINPUT95), .B2(new_n265), .ZN(new_n269));
  OR2_X1    g068(.A1(G71gat), .A2(G78gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n270), .B1(KEYINPUT94), .B2(new_n267), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(KEYINPUT94), .B2(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n267), .B1(new_n270), .B2(new_n266), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n269), .A2(new_n272), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT21), .ZN(new_n275));
  AND2_X1   g074(.A1(G231gat), .A2(G233gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G127gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G15gat), .B(G22gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT16), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(G1gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT91), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n281), .B(new_n282), .C1(G1gat), .C2(new_n279), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n283), .A2(G8gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(G8gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n286), .B1(KEYINPUT21), .B2(new_n274), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n278), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G183gat), .B(G211gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n289), .B(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n202), .B1(new_n264), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n294), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n289), .B(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n298), .A2(new_n259), .A3(KEYINPUT99), .A4(new_n263), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G230gat), .ZN(new_n301));
  INV_X1    g100(.A(G233gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT10), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n269), .A2(new_n272), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n273), .A2(new_n265), .ZN(new_n306));
  INV_X1    g105(.A(new_n235), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(new_n306), .C1(new_n233), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n274), .B1(new_n236), .B2(new_n238), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n304), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n242), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n303), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n303), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OR3_X1    g118(.A1(new_n313), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n313), .B2(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n300), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT72), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n252), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g128(.A1(G211gat), .A2(G218gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G197gat), .ZN(new_n333));
  INV_X1    g132(.A(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n335), .A2(new_n336), .B1(new_n338), .B2(new_n330), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n326), .A3(new_n331), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(KEYINPUT73), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT73), .B1(new_n341), .B2(new_n343), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT23), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n354), .A2(new_n355), .A3(new_n360), .A4(KEYINPUT25), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT25), .A4(new_n353), .ZN(new_n362));
  AND2_X1   g161(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n357), .A2(new_n356), .B1(new_n363), .B2(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT66), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n358), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n368), .A2(new_n369), .B1(new_n357), .B2(new_n356), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT65), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n375), .A3(new_n354), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G226gat), .A2(G233gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n348), .A2(new_n349), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n353), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT26), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n357), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT28), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G183gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT67), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n241), .ZN(new_n390));
  INV_X1    g189(.A(G183gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT27), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n388), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n385), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n385), .A2(G190gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n387), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT68), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n395), .A2(new_n387), .A3(new_n392), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n384), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n378), .A2(new_n379), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n379), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n354), .B1(new_n374), .B2(KEYINPUT65), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n370), .A2(KEYINPUT65), .A3(new_n358), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n377), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n361), .A2(new_n365), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n401), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n404), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n347), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n409), .A2(G226gat), .A3(new_n410), .A4(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n414));
  INV_X1    g213(.A(new_n343), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n342), .B1(new_n326), .B2(new_n331), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n344), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n378), .A2(new_n401), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n413), .B(new_n418), .C1(new_n419), .C2(new_n404), .ZN(new_n420));
  XOR2_X1   g219(.A(G8gat), .B(G36gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT74), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n412), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n412), .B2(new_n420), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT30), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n428), .B(new_n424), .C1(new_n412), .C2(new_n420), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G120gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G113gat), .ZN(new_n432));
  INV_X1    g231(.A(G113gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G120gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT69), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n437));
  INV_X1    g236(.A(G134gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G127gat), .ZN(new_n439));
  INV_X1    g238(.A(G127gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G134gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n437), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT1), .B1(new_n432), .B2(new_n434), .ZN(new_n444));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n436), .A2(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT70), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n439), .A2(new_n441), .ZN(new_n448));
  XNOR2_X1  g247(.A(G113gat), .B(G120gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(KEYINPUT1), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n450), .B(new_n451), .C1(new_n436), .C2(new_n443), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G141gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G148gat), .ZN(new_n456));
  INV_X1    g255(.A(G148gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G141gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G155gat), .B(G162gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT2), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT77), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n456), .A2(new_n458), .B1(KEYINPUT2), .B2(new_n461), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n462), .ZN(new_n468));
  INV_X1    g267(.A(new_n461), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT75), .ZN(new_n470));
  INV_X1    g269(.A(G162gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n291), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n474), .B2(KEYINPUT76), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476));
  AOI211_X1 g275(.A(new_n476), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n464), .B(new_n467), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT80), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n454), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  AND4_X1   g281(.A1(new_n466), .A2(new_n459), .A3(new_n460), .A4(new_n462), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n466), .B1(new_n465), .B2(new_n460), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n473), .ZN(new_n486));
  NOR3_X1   g285(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n461), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n476), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT76), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n468), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n485), .A2(new_n447), .A3(new_n491), .A4(new_n452), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT80), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g292(.A(new_n446), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n481), .B1(new_n479), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n482), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n478), .B2(KEYINPUT3), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n485), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT81), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n502), .ZN(new_n505));
  AOI211_X1 g304(.A(KEYINPUT5), .B(new_n505), .C1(new_n497), .C2(new_n499), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT81), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n485), .A2(new_n491), .A3(new_n494), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(KEYINPUT80), .C1(KEYINPUT4), .C2(new_n492), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n506), .A2(new_n507), .A3(new_n510), .A4(new_n482), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n446), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT78), .A3(new_n508), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n478), .A2(new_n514), .A3(new_n446), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n505), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n454), .A2(KEYINPUT4), .A3(new_n479), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n481), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n500), .A2(new_n518), .A3(new_n502), .A4(new_n519), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n504), .A2(new_n511), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G1gat), .B(G29gat), .Z(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G57gat), .B(G85gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT6), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n511), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n517), .A2(new_n520), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(KEYINPUT6), .A3(new_n531), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n430), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT83), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G228gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n341), .A2(new_n403), .A3(new_n343), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT82), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n341), .A2(new_n543), .A3(new_n403), .A4(new_n343), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n498), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n478), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n403), .B1(new_n478), .B2(KEYINPUT3), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n347), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n540), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n418), .B1(new_n403), .B2(new_n499), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n415), .A2(new_n416), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n478), .A2(new_n551), .A3(new_n403), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n478), .A2(KEYINPUT3), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n540), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G78gat), .B(G106gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT31), .B(G50gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  NOR3_X1   g357(.A1(new_n549), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT3), .B1(new_n541), .B2(KEYINPUT82), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n479), .B1(new_n561), .B2(new_n544), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n539), .B1(new_n550), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n553), .A3(new_n540), .A4(new_n552), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n538), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n558), .B1(new_n549), .B2(new_n555), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n563), .A2(new_n564), .A3(new_n560), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n537), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT84), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G15gat), .B(G43gat), .Z(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G99gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G227gat), .A2(G233gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n453), .B1(new_n378), .B2(new_n401), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n409), .A2(new_n454), .A3(new_n410), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n579), .B2(KEYINPUT33), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n578), .ZN(new_n584));
  INV_X1    g383(.A(new_n576), .ZN(new_n585));
  AOI221_X4 g384(.A(new_n581), .B1(KEYINPUT33), .B2(new_n575), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT71), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n577), .A2(new_n576), .A3(new_n578), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT34), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n378), .A2(new_n453), .A3(new_n401), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n454), .B1(new_n409), .B2(new_n410), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n595), .A3(new_n575), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n582), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n587), .A2(new_n589), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n588), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(KEYINPUT36), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n589), .B1(new_n583), .B2(new_n586), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n583), .A2(new_n589), .A3(new_n586), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n536), .A2(new_n572), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n521), .A2(new_n611), .A3(new_n526), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT88), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n526), .B(KEYINPUT85), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n530), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT88), .A2(new_n612), .B1(new_n527), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n412), .A2(new_n420), .A3(KEYINPUT37), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT38), .B1(new_n618), .B2(KEYINPUT87), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n424), .A2(KEYINPUT37), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n425), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n619), .B(new_n621), .C1(KEYINPUT87), .C2(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT38), .ZN(new_n624));
  INV_X1    g423(.A(new_n426), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n617), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n530), .A2(new_n615), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n427), .A2(new_n429), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n482), .B(new_n500), .C1(new_n493), .C2(new_n495), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n505), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT86), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n631), .A2(KEYINPUT86), .A3(new_n505), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n615), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n513), .A2(new_n515), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(new_n502), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n639), .B1(new_n638), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n630), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n569), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n537), .B1(new_n567), .B2(new_n568), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n627), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n528), .A2(new_n526), .A3(new_n529), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n611), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n521), .A2(new_n526), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n534), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n608), .A2(new_n570), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n653), .A2(new_n629), .A3(new_n654), .A4(new_n600), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT35), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n427), .A2(KEYINPUT35), .A3(new_n429), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(new_n606), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT88), .ZN(new_n659));
  OAI22_X1  g458(.A1(new_n628), .A2(new_n651), .B1(new_n534), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n654), .B(new_n658), .C1(new_n660), .C2(new_n613), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n610), .A2(new_n649), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT18), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT92), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n286), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n223), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n243), .A2(new_n286), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(KEYINPUT93), .B(new_n663), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n286), .B(new_n243), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n669), .B(KEYINPUT13), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n666), .A2(new_n669), .A3(new_n667), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n333), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT11), .B(G169gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT12), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n682), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n671), .A2(new_n684), .A3(new_n674), .A4(new_n676), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n323), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n653), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g492(.A1(new_n689), .A2(new_n629), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT101), .ZN(new_n697));
  OAI21_X1  g496(.A(G8gat), .B1(new_n689), .B2(new_n629), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n697), .B(new_n699), .C1(KEYINPUT42), .C2(new_n700), .ZN(G1325gat));
  NOR2_X1   g500(.A1(new_n607), .A2(new_n608), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n689), .A2(G15gat), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n604), .A2(new_n609), .ZN(new_n705));
  OAI21_X1  g504(.A(G15gat), .B1(new_n689), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n572), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT103), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(new_n264), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n662), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n322), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n295), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n687), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(G29gat), .A3(new_n653), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT45), .Z(new_n720));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT35), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n603), .A2(new_n569), .A3(new_n566), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n596), .A2(new_n597), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n602), .B1(new_n724), .B2(KEYINPUT71), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n599), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n722), .B1(new_n726), .B2(new_n535), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n657), .A2(new_n648), .A3(new_n603), .A4(new_n606), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n614), .B2(new_n617), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n721), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n656), .A2(KEYINPUT104), .A3(new_n661), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(new_n731), .B1(new_n649), .B2(new_n610), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n610), .A2(new_n649), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n727), .A2(new_n729), .A3(new_n721), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT104), .B1(new_n656), .B2(new_n661), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n733), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n662), .B2(new_n713), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n735), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n717), .ZN(new_n744));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744), .B2(new_n653), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n720), .A2(new_n745), .ZN(G1328gat));
  OR3_X1    g545(.A1(new_n718), .A2(G36gat), .A3(new_n629), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G36gat), .B1(new_n744), .B2(new_n629), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(KEYINPUT46), .A3(new_n749), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(G1329gat));
  INV_X1    g554(.A(new_n705), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n743), .A2(new_n756), .A3(new_n717), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n718), .A2(G43gat), .A3(new_n703), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT107), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT107), .B(new_n762), .C1(new_n758), .C2(new_n759), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(G1330gat));
  OAI21_X1  g563(.A(G50gat), .B1(new_n744), .B2(new_n648), .ZN(new_n765));
  INV_X1    g564(.A(new_n572), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n713), .A2(new_n716), .A3(G50gat), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n688), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n688), .A2(new_n767), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n743), .A2(new_n572), .A3(new_n717), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g572(.A1(new_n732), .A2(new_n300), .A3(new_n686), .A4(new_n715), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n691), .ZN(new_n775));
  XNOR2_X1  g574(.A(KEYINPUT108), .B(G57gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1332gat));
  AOI21_X1  g576(.A(new_n629), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n779), .B(new_n780), .Z(G1333gat));
  INV_X1    g580(.A(G71gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n774), .A2(new_n782), .A3(new_n702), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n774), .A2(new_n756), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n572), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g587(.A1(new_n295), .A2(new_n687), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n715), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n743), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n743), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n653), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n713), .A2(new_n789), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n739), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n691), .A2(new_n230), .A3(new_n322), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n796), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  OAI21_X1  g604(.A(KEYINPUT112), .B1(new_n791), .B2(new_n629), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n743), .A2(new_n807), .A3(new_n430), .A4(new_n790), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(G92gat), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n430), .A2(new_n322), .A3(new_n231), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT110), .Z(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n800), .B2(new_n801), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT111), .B(new_n812), .C1(new_n800), .C2(new_n801), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n792), .A2(new_n430), .A3(new_n794), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n813), .B1(new_n819), .B2(G92gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n810), .ZN(G1337gat));
  OAI21_X1  g620(.A(G99gat), .B1(new_n795), .B2(new_n705), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n703), .A2(G99gat), .A3(new_n715), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT113), .Z(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n803), .B2(new_n824), .ZN(G1338gat));
  OAI21_X1  g624(.A(G106gat), .B1(new_n791), .B2(new_n648), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n715), .A2(G106gat), .A3(new_n648), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT53), .B1(new_n802), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n827), .B(KEYINPUT114), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n803), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n792), .A2(new_n572), .A3(new_n794), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n833), .B2(new_n834), .ZN(G1339gat));
  AOI21_X1  g634(.A(new_n669), .B1(new_n666), .B2(new_n667), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n672), .A2(new_n673), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n681), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n685), .A2(new_n322), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n318), .B1(new_n313), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n274), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n242), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT10), .B1(new_n843), .B2(new_n308), .ZN(new_n844));
  INV_X1    g643(.A(new_n312), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n314), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n311), .A2(new_n303), .A3(new_n312), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT54), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n841), .A2(new_n848), .A3(new_n849), .A4(KEYINPUT55), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n320), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n841), .A2(new_n848), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n686), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n264), .B1(new_n839), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n685), .A2(new_n838), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n858), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n263), .B2(new_n259), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n295), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n296), .A2(new_n299), .A3(new_n687), .A4(new_n715), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n653), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n629), .A3(new_n726), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT117), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n433), .A3(new_n686), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n572), .B(new_n703), .C1(new_n861), .C2(new_n862), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n691), .A2(new_n629), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n871), .A2(new_n686), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n866), .B1(new_n873), .B2(new_n433), .ZN(G1340gat));
  NAND2_X1  g673(.A1(new_n322), .A2(new_n431), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT118), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n871), .A2(new_n322), .A3(new_n872), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n431), .ZN(G1341gat));
  AND3_X1   g678(.A1(new_n871), .A2(new_n298), .A3(new_n872), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n298), .A2(new_n440), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n880), .A2(new_n440), .B1(new_n864), .B2(new_n881), .ZN(G1342gat));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n438), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n864), .A2(new_n713), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n871), .A2(new_n264), .A3(new_n872), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n438), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n869), .A2(new_n705), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n648), .B1(new_n861), .B2(new_n862), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n855), .A2(new_n320), .A3(new_n850), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n841), .A2(new_n848), .A3(KEYINPUT121), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT121), .B1(new_n841), .B2(new_n848), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n897), .A2(KEYINPUT55), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT122), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(KEYINPUT55), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n896), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n902), .A2(new_n851), .A3(new_n903), .A4(new_n855), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n686), .A3(new_n904), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n839), .B(KEYINPUT120), .Z(new_n906));
  AOI21_X1  g705(.A(new_n264), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n295), .B1(new_n907), .B2(new_n860), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n766), .B1(new_n908), .B2(new_n862), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n894), .B1(new_n893), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n687), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n863), .A2(new_n629), .A3(new_n570), .A4(new_n705), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n455), .A3(new_n686), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT58), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1344gat));
  NAND3_X1  g718(.A1(new_n913), .A2(new_n457), .A3(new_n322), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n910), .A2(new_n715), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(KEYINPUT59), .A3(new_n457), .ZN(new_n922));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n862), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n893), .A3(new_n572), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n861), .A2(new_n862), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT57), .B1(new_n926), .B2(new_n648), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n715), .B1(new_n891), .B2(KEYINPUT124), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n923), .B1(new_n930), .B2(G148gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n920), .B1(new_n922), .B2(new_n931), .ZN(G1345gat));
  OAI21_X1  g731(.A(G155gat), .B1(new_n910), .B2(new_n295), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n291), .A3(new_n298), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1346gat));
  NOR3_X1   g734(.A1(new_n910), .A2(new_n471), .A3(new_n713), .ZN(new_n936));
  AOI21_X1  g735(.A(G162gat), .B1(new_n913), .B2(new_n264), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  AOI21_X1  g737(.A(new_n691), .B1(new_n861), .B2(new_n862), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n726), .A2(new_n430), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT125), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n348), .A3(new_n686), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n691), .A2(new_n629), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n867), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n686), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT126), .A3(G169gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT126), .B1(new_n948), .B2(G169gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(G1348gat));
  OAI21_X1  g750(.A(G176gat), .B1(new_n946), .B2(new_n715), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n943), .A2(new_n349), .A3(new_n322), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  OAI21_X1  g753(.A(G183gat), .B1(new_n946), .B2(new_n295), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n298), .A2(new_n387), .A3(new_n392), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n942), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n241), .A3(new_n264), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n947), .A2(new_n264), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(G190gat), .ZN(new_n962));
  AOI211_X1 g761(.A(KEYINPUT61), .B(new_n241), .C1(new_n947), .C2(new_n264), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(G1351gat));
  AND2_X1   g763(.A1(new_n945), .A2(new_n705), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n925), .A2(new_n927), .A3(new_n965), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(new_n333), .A3(new_n687), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n756), .A2(new_n629), .A3(new_n648), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n939), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n686), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n967), .A2(new_n971), .ZN(G1352gat));
  NAND4_X1  g771(.A1(new_n925), .A2(new_n927), .A3(new_n322), .A4(new_n965), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G204gat), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n715), .A2(G204gat), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(KEYINPUT62), .B1(new_n969), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n939), .A2(new_n978), .A3(new_n968), .A4(new_n975), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n974), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n327), .A3(new_n298), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n925), .A2(new_n927), .A3(new_n298), .A4(new_n965), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n987), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n987), .B2(G211gat), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(G1354gat));
  OAI21_X1  g789(.A(G218gat), .B1(new_n966), .B2(new_n713), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n252), .A3(new_n264), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1355gat));
endmodule


