//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT96), .B1(new_n202), .B2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G22gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G15gat), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(G8gat), .B1(new_n203), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n207), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(new_n208), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n214), .A2(KEYINPUT96), .A3(new_n215), .A4(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G43gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G50gat), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT15), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT92), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G29gat), .A2(G36gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n222), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT94), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(new_n218), .B2(G50gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n220), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n219), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n223), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n222), .A3(new_n232), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n241), .A2(new_n222), .A3(new_n232), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n239), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT94), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n233), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n217), .B1(new_n247), .B2(KEYINPUT17), .ZN(new_n248));
  INV_X1    g047(.A(new_n233), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n240), .A2(new_n242), .A3(new_n234), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT94), .B1(new_n244), .B2(new_n245), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT95), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n247), .A2(new_n255), .A3(KEYINPUT17), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n248), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT98), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n212), .A2(KEYINPUT97), .A3(new_n216), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT97), .B1(new_n212), .B2(new_n216), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n247), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT97), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n217), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n212), .A2(KEYINPUT97), .A3(new_n216), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT98), .A3(new_n252), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G229gat), .A2(G233gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n257), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT18), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n257), .A2(new_n268), .A3(KEYINPUT18), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n247), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n269), .B(KEYINPUT13), .Z(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G141gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G169gat), .B(G197gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT12), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n272), .A2(new_n273), .A3(new_n277), .A4(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G1gat), .B(G29gat), .Z(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G57gat), .B(G85gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G127gat), .B(G134gat), .Z(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n296), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(KEYINPUT1), .ZN(new_n302));
  INV_X1    g101(.A(G113gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G120gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT70), .B(G120gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310));
  XNOR2_X1  g109(.A(G155gat), .B(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT79), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315));
  AND2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT80), .B(G162gat), .Z(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n314), .A3(new_n311), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n309), .A2(new_n310), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT84), .B1(new_n324), .B2(new_n308), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n323), .A2(new_n325), .B1(new_n324), .B2(new_n308), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n318), .A2(new_n322), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n309), .B1(KEYINPUT3), .B2(new_n324), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n323), .A2(new_n325), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n324), .B(KEYINPUT83), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT85), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT85), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n335), .A2(new_n343), .A3(new_n338), .A4(new_n340), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n328), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n337), .A3(new_n309), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n337), .B1(new_n323), .B2(new_n325), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT87), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n347), .ZN(new_n353));
  AOI211_X1 g152(.A(KEYINPUT5), .B(new_n329), .C1(new_n333), .C2(new_n334), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n294), .B1(new_n346), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n333), .A2(new_n334), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n350), .A2(new_n357), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n329), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT39), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n326), .B2(new_n327), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n360), .A3(new_n329), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n294), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT40), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n356), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G8gat), .B(G36gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  INV_X1    g168(.A(G226gat), .ZN(new_n370));
  INV_X1    g169(.A(G233gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT23), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT25), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n374), .B2(KEYINPUT23), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n382), .B(KEYINPUT67), .Z(new_n383));
  INV_X1    g182(.A(KEYINPUT24), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(G183gat), .A3(G190gat), .ZN(new_n385));
  AND2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n384), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n382), .B(KEYINPUT64), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT65), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(KEYINPUT65), .A3(new_n387), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT66), .B1(new_n375), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n396), .A3(KEYINPUT23), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n395), .A2(new_n397), .B1(new_n375), .B2(new_n377), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n388), .B1(new_n399), .B2(new_n379), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT27), .B(G183gat), .ZN(new_n401));
  INV_X1    g200(.A(G190gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n403), .A2(KEYINPUT68), .A3(KEYINPUT28), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n402), .B2(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n375), .A2(new_n407), .A3(new_n376), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n386), .B1(KEYINPUT26), .B2(new_n374), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n404), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n373), .B1(new_n412), .B2(KEYINPUT29), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT73), .B(G218gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT22), .B1(new_n414), .B2(G211gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT74), .ZN(new_n416));
  XNOR2_X1  g215(.A(G197gat), .B(G204gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n379), .ZN(new_n424));
  INV_X1    g223(.A(new_n388), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n411), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT76), .B1(new_n428), .B2(new_n372), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n412), .A2(new_n430), .A3(new_n373), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n413), .B(new_n423), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n372), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n423), .B(KEYINPUT75), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n369), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT77), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(new_n369), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT78), .A4(new_n369), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT30), .A4(new_n369), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n438), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n362), .A2(KEYINPUT40), .A3(new_n294), .A4(new_n363), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n366), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n442), .A2(new_n444), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT90), .ZN(new_n451));
  OR3_X1    g250(.A1(new_n434), .A2(new_n435), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n434), .B2(new_n435), .ZN(new_n453));
  INV_X1    g252(.A(new_n423), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n429), .A2(new_n431), .ZN(new_n455));
  INV_X1    g254(.A(new_n413), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT38), .B1(new_n458), .B2(KEYINPUT37), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n369), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n437), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n450), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n346), .A2(new_n294), .A3(new_n355), .ZN(new_n465));
  INV_X1    g264(.A(new_n294), .ZN(new_n466));
  INV_X1    g265(.A(new_n355), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n345), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n356), .A2(new_n469), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n460), .B1(new_n432), .B2(new_n436), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT38), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n464), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G228gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n371), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n324), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT29), .B1(new_n421), .B2(new_n422), .ZN(new_n480));
  INV_X1    g279(.A(new_n330), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT29), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n333), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n482), .A2(new_n483), .B1(new_n454), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(KEYINPUT89), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n477), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n480), .A2(new_n324), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n477), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n435), .B2(new_n485), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n488), .A2(G22gat), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n482), .A2(new_n483), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n485), .A2(new_n454), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n487), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n477), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n435), .A2(new_n485), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n490), .A3(new_n477), .A4(new_n489), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n204), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(G78gat), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(G22gat), .B1(new_n488), .B2(new_n492), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n500), .A3(new_n204), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT31), .B(G50gat), .ZN(new_n507));
  INV_X1    g306(.A(G106gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n502), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n503), .B2(new_n504), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n449), .A2(new_n475), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n471), .A2(new_n472), .ZN(new_n516));
  INV_X1    g315(.A(new_n447), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n426), .A2(new_n308), .A3(new_n427), .ZN(new_n523));
  AND2_X1   g322(.A1(G227gat), .A2(G233gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n309), .B1(new_n400), .B2(new_n411), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT32), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G43gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n526), .B(KEYINPUT32), .C1(new_n534), .C2(new_n533), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n523), .A2(new_n525), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(new_n524), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n522), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n539), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n537), .A3(new_n540), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n521), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n547), .A3(KEYINPUT36), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n547), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n515), .A2(new_n520), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n514), .A2(new_n510), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT35), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n447), .B1(new_n472), .B2(new_n471), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n549), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n514), .A2(new_n510), .A3(new_n549), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT35), .B1(new_n557), .B2(new_n518), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n289), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n516), .ZN(new_n561));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g362(.A(G71gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n505), .ZN(new_n565));
  XNOR2_X1  g364(.A(G57gat), .B(G64gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G64gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G57gat), .ZN(new_n570));
  INV_X1    g369(.A(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G64gat), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n570), .A2(new_n572), .A3(new_n567), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n562), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT100), .B(G57gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n575), .B2(new_n569), .ZN(new_n576));
  INV_X1    g375(.A(new_n562), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n577), .A3(new_n565), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n266), .B1(KEYINPUT21), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT102), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G155gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT101), .B(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G127gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n592), .B(new_n593), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n586), .A3(new_n585), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT104), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT8), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n603), .A2(new_n606), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n606), .A4(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  OR3_X1    g417(.A1(new_n611), .A2(new_n614), .A3(new_n612), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n252), .B2(new_n253), .ZN(new_n621));
  INV_X1    g420(.A(new_n254), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n252), .A2(KEYINPUT95), .A3(new_n253), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n618), .A2(new_n619), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n252), .A2(new_n625), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n601), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n601), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n254), .A2(new_n256), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n631), .B(new_n628), .C1(new_n632), .C2(new_n621), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n630), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n630), .B2(new_n633), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n599), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n625), .A2(new_n579), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n613), .A2(new_n617), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n574), .A2(new_n647), .A3(new_n578), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT10), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n620), .A2(new_n650), .A3(new_n579), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT105), .ZN(new_n653));
  INV_X1    g452(.A(new_n645), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n618), .A2(new_n619), .B1(new_n574), .B2(new_n578), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n574), .A2(new_n647), .A3(new_n578), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n580), .A2(new_n625), .A3(KEYINPUT10), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n655), .A2(new_n656), .A3(new_n645), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n644), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n659), .A2(new_n663), .A3(new_n644), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n640), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n560), .A2(new_n561), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT106), .B(G1gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  NAND3_X1  g472(.A1(new_n560), .A2(new_n447), .A3(new_n670), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT16), .B(G8gat), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT107), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(G8gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(G1325gat));
  NAND4_X1  g479(.A1(new_n560), .A2(new_n206), .A3(new_n549), .A4(new_n670), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n560), .A2(new_n670), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n543), .A2(new_n547), .A3(KEYINPUT36), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT36), .B1(new_n543), .B2(new_n547), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT108), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n551), .A2(new_n687), .A3(new_n548), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n682), .B1(new_n690), .B2(G15gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT109), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n683), .A2(new_n519), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT43), .B(G22gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NAND2_X1  g494(.A1(new_n552), .A2(new_n559), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n599), .A2(new_n668), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n289), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n696), .A2(new_n639), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n228), .A3(new_n561), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n639), .ZN(new_n702));
  INV_X1    g501(.A(new_n639), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n515), .A2(new_n520), .A3(new_n686), .A4(new_n688), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n559), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n702), .B(new_n698), .C1(KEYINPUT44), .C2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n516), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n707), .ZN(G1328gat));
  NOR2_X1   g507(.A1(new_n517), .A2(G36gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT110), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n699), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n706), .B2(new_n517), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT46), .B1(new_n711), .B2(new_n713), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  NAND2_X1  g517(.A1(new_n689), .A2(G43gat), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n706), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n697), .A2(new_n703), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n560), .A2(new_n549), .A3(new_n723), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n724), .A2(new_n218), .B1(new_n721), .B2(KEYINPUT47), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n722), .B1(new_n720), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(G1330gat));
  OAI21_X1  g527(.A(G50gat), .B1(new_n706), .B2(new_n553), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT48), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n699), .A2(new_n220), .A3(new_n519), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n729), .B(new_n732), .C1(new_n730), .C2(KEYINPUT48), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1331gat));
  NAND3_X1  g535(.A1(new_n640), .A2(new_n289), .A3(new_n667), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n559), .B2(new_n704), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n561), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n575), .ZN(G1332gat));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n447), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT49), .B(G64gat), .Z(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n741), .B2(new_n743), .ZN(G1333gat));
  AOI21_X1  g543(.A(new_n564), .B1(new_n738), .B2(new_n689), .ZN(new_n745));
  INV_X1    g544(.A(new_n549), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(G71gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n738), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n519), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  INV_X1    g551(.A(new_n599), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(new_n288), .A3(new_n668), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n702), .B(new_n754), .C1(KEYINPUT44), .C2(new_n705), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n516), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n668), .A2(G85gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n561), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n753), .A2(new_n288), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT51), .B1(new_n705), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n760), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n752), .B1(new_n757), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n764), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(KEYINPUT113), .A3(new_n756), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1336gat));
  OAI21_X1  g567(.A(G92gat), .B1(new_n755), .B2(new_n517), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n517), .A2(G92gat), .A3(new_n668), .ZN(new_n771));
  INV_X1    g570(.A(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n772), .B2(new_n761), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n774), .A3(KEYINPUT52), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n769), .B(new_n773), .C1(KEYINPUT114), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1337gat));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT115), .B(G99gat), .Z(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n549), .A3(new_n667), .A4(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n689), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n755), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n783), .B2(new_n780), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n755), .B2(new_n553), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n668), .A2(G106gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n519), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n762), .B2(new_n763), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n789), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n792), .A3(new_n785), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1339gat));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n657), .A2(new_n658), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n645), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n657), .A2(new_n654), .A3(new_n658), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n653), .A2(new_n661), .A3(new_n796), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n801), .A3(new_n644), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT116), .A4(new_n644), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n799), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n801), .A2(new_n644), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n665), .B1(new_n808), .B2(new_n795), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n288), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n257), .A2(new_n268), .ZN(new_n811));
  INV_X1    g610(.A(new_n269), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n276), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n268), .A2(new_n274), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n816), .A2(new_n817), .A3(new_n283), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n816), .B2(new_n283), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n667), .B(new_n287), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n639), .B1(new_n810), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n639), .B(new_n287), .C1(new_n818), .C2(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n809), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n599), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n640), .A2(new_n289), .A3(new_n668), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n516), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n557), .A2(new_n447), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n288), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n519), .B1(new_n825), .B2(new_n826), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n746), .A2(new_n516), .A3(new_n447), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(new_n303), .A3(new_n289), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n830), .A2(new_n834), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n833), .B2(new_n668), .ZN(new_n836));
  INV_X1    g635(.A(new_n829), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n668), .A2(new_n305), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G1341gat));
  OAI21_X1  g638(.A(G127gat), .B1(new_n833), .B2(new_n599), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n599), .A2(G127gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n837), .B2(new_n841), .ZN(G1342gat));
  OR3_X1    g641(.A1(new_n837), .A2(G134gat), .A3(new_n703), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT118), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n831), .A2(new_n639), .A3(new_n832), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n846), .B2(G134gat), .ZN(new_n847));
  INV_X1    g646(.A(new_n843), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n782), .A2(new_n519), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n827), .A2(new_n517), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n782), .A2(KEYINPUT121), .A3(new_n519), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n289), .A2(G141gat), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT58), .B1(new_n856), .B2(KEYINPUT122), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n825), .A2(new_n826), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n519), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n516), .A2(new_n447), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n782), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n820), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n289), .B1(new_n823), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n806), .A2(KEYINPUT119), .A3(new_n809), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n639), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n599), .B1(new_n869), .B2(new_n824), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n553), .B1(new_n870), .B2(new_n826), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n871), .B2(new_n860), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT123), .B1(new_n872), .B2(new_n289), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G141gat), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(KEYINPUT123), .A3(new_n289), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n857), .B(new_n858), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n856), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n863), .B(KEYINPUT120), .C1(new_n871), .C2(new_n860), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n288), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n877), .B1(new_n881), .B2(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(G1344gat));
  NAND3_X1  g683(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(G148gat), .A3(new_n668), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n860), .B1(new_n859), .B2(new_n519), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n887), .B1(new_n871), .B2(new_n860), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n667), .A3(new_n782), .A4(new_n862), .ZN(new_n889));
  AND2_X1   g688(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n879), .A2(new_n880), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n894), .B2(new_n667), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n891), .B1(new_n895), .B2(KEYINPUT59), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n893), .B2(new_n599), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n753), .A2(new_n320), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n885), .B2(new_n898), .ZN(G1346gat));
  NOR2_X1   g698(.A1(new_n893), .A2(new_n703), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n639), .A2(new_n319), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n900), .A2(new_n319), .B1(new_n885), .B2(new_n901), .ZN(G1347gat));
  NAND4_X1  g701(.A1(new_n831), .A2(new_n516), .A3(new_n447), .A4(new_n549), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n289), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n859), .B2(new_n516), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT124), .B(new_n561), .C1(new_n825), .C2(new_n826), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n557), .A2(new_n517), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n288), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n913), .B2(new_n904), .ZN(G1348gat));
  OAI21_X1  g713(.A(G176gat), .B1(new_n903), .B2(new_n668), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n668), .A2(G176gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n911), .B2(new_n916), .ZN(G1349gat));
  OAI21_X1  g716(.A(G183gat), .B1(new_n903), .B2(new_n599), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n753), .A2(new_n401), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n912), .A2(new_n402), .A3(new_n639), .ZN(new_n922));
  OAI21_X1  g721(.A(G190gat), .B1(new_n903), .B2(new_n703), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n689), .A2(new_n561), .A3(new_n517), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n888), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(G197gat), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n927), .A2(new_n928), .A3(new_n289), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n447), .A2(new_n686), .A3(new_n688), .A4(new_n519), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n907), .B2(new_n908), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT125), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n930), .B(new_n933), .C1(new_n907), .C2(new_n908), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n288), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n929), .B1(new_n928), .B2(new_n935), .ZN(G1352gat));
  OR3_X1    g735(.A1(new_n931), .A2(G204gat), .A3(new_n668), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n927), .B2(new_n668), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G1353gat));
  NOR2_X1   g740(.A1(new_n599), .A2(G211gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n932), .A2(new_n934), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n888), .A2(new_n753), .A3(new_n926), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  NAND4_X1  g746(.A1(new_n888), .A2(new_n414), .A3(new_n639), .A4(new_n926), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n639), .A3(new_n934), .ZN(new_n949));
  INV_X1    g748(.A(G218gat), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n949), .A2(KEYINPUT126), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT126), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n948), .C1(new_n951), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1355gat));
endmodule


