//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n207), .A2(G169gat), .A3(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n204), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT27), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT69), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n219), .A2(KEYINPUT28), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(G190gat), .B1(new_n212), .B2(KEYINPUT68), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT28), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n202), .B(new_n210), .C1(new_n221), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n202), .A2(KEYINPUT24), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(G183gat), .A3(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n203), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n232), .A2(new_n234), .B1(new_n206), .B2(new_n208), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n237));
  OAI21_X1  g036(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n238));
  OR3_X1    g037(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n240), .B2(new_n235), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n236), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI211_X1 g042(.A(KEYINPUT67), .B(new_n237), .C1(new_n240), .C2(new_n235), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n226), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G134gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G127gat), .ZN(new_n247));
  INV_X1    g046(.A(G127gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G134gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT70), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251));
  OAI221_X1 g050(.A(new_n250), .B1(KEYINPUT70), .B2(new_n247), .C1(KEYINPUT1), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253));
  INV_X1    g052(.A(G113gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(G120gat), .A3(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n254), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(KEYINPUT72), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n247), .A2(new_n249), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT72), .B1(new_n257), .B2(new_n259), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n226), .B(new_n265), .C1(new_n243), .C2(new_n244), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G227gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT34), .ZN(new_n274));
  AOI22_X1  g073(.A1(new_n269), .A2(new_n273), .B1(KEYINPUT74), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n267), .A2(new_n272), .A3(new_n268), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n280));
  XOR2_X1   g079(.A(G71gat), .B(G99gat), .Z(new_n281));
  XNOR2_X1  g080(.A(G15gat), .B(G43gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n280), .B1(new_n283), .B2(KEYINPUT33), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(KEYINPUT33), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(KEYINPUT73), .A2(new_n285), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n289), .A3(new_n284), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n278), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n283), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(KEYINPUT73), .ZN(new_n293));
  AND4_X1   g092(.A1(new_n278), .A2(new_n292), .A3(new_n293), .A4(new_n290), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n276), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n290), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n277), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(new_n278), .A3(new_n290), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n298), .A3(new_n275), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(KEYINPUT36), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n297), .A2(new_n298), .A3(new_n275), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n275), .B1(new_n297), .B2(new_n298), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G8gat), .B(G36gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G64gat), .B(G92gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n245), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n226), .B(new_n310), .C1(new_n243), .C2(new_n244), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(KEYINPUT22), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(new_n322), .A3(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n308), .B1(new_n326), .B2(KEYINPUT37), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT37), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT38), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n325), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n322), .B1(new_n313), .B2(new_n314), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n308), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n308), .A2(KEYINPUT37), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n328), .B1(new_n331), .B2(KEYINPUT84), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n324), .A2(new_n337), .A3(new_n325), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT38), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n307), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n330), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n344), .ZN(new_n350));
  AND2_X1   g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n344), .A2(new_n354), .A3(KEYINPUT2), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n346), .A2(new_n350), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n345), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  AND2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT4), .B1(new_n265), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n257), .A2(new_n259), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(new_n260), .A3(new_n262), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n356), .A2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .A4(new_n252), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n356), .A2(new_n365), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n377), .B1(new_n356), .B2(new_n365), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n265), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n375), .A2(new_n376), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n265), .A2(new_n366), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(new_n372), .A3(new_n252), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n376), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n383), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT78), .B(KEYINPUT0), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT79), .ZN(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n394), .B(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n398), .A3(new_n388), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n367), .A2(new_n374), .B1(new_n265), .B2(new_n380), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n383), .A3(new_n376), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n390), .A2(new_n397), .A3(new_n399), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n390), .A2(new_n399), .A3(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n397), .B1(new_n405), .B2(KEYINPUT83), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n390), .A2(new_n407), .A3(new_n399), .A4(new_n401), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n394), .B(new_n395), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n343), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n322), .A2(new_n311), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n372), .B1(new_n414), .B2(new_n377), .ZN(new_n415));
  INV_X1    g214(.A(new_n378), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n322), .B1(new_n416), .B2(new_n311), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n417), .A2(new_n421), .B1(new_n422), .B2(new_n271), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G22gat), .ZN(new_n424));
  INV_X1    g223(.A(G22gat), .ZN(new_n425));
  OAI221_X1 g224(.A(new_n425), .B1(new_n422), .B2(new_n271), .C1(new_n417), .C2(new_n421), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT31), .B(G50gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n424), .B2(new_n426), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n420), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n424), .A2(new_n426), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n427), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n429), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n405), .A2(KEYINPUT83), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n410), .A3(new_n408), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n324), .A2(KEYINPUT30), .A3(new_n325), .A4(new_n307), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n333), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n342), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n400), .A2(KEYINPUT39), .A3(new_n376), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT82), .B1(new_n447), .B2(new_n410), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n375), .A2(new_n381), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n387), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n397), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n400), .A2(new_n376), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT39), .B1(new_n386), .B2(new_n387), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n446), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  AOI211_X1 g258(.A(KEYINPUT40), .B(new_n457), .C1(new_n448), .C2(new_n453), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n437), .B1(new_n445), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n300), .B(new_n304), .C1(new_n413), .C2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT81), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT81), .B1(new_n432), .B2(new_n436), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n405), .A2(new_n410), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n403), .A3(new_n402), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n444), .B1(new_n468), .B2(new_n411), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  INV_X1    g270(.A(new_n437), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n295), .B2(new_n299), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n473), .B2(new_n469), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n437), .B1(new_n302), .B2(new_n303), .ZN(new_n475));
  INV_X1    g274(.A(new_n444), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n471), .B(new_n476), .C1(new_n409), .C2(new_n412), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI22_X1  g277(.A1(new_n463), .A2(new_n470), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT18), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  INV_X1    g281(.A(G29gat), .ZN(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT14), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(G29gat), .B2(G36gat), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT86), .B(G36gat), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(G29gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(new_n487), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n494), .A2(new_n495), .B1(new_n490), .B2(G29gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n482), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT17), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(G1gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT16), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n503), .B2(G1gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n502), .B(new_n504), .C1(new_n506), .C2(G8gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n493), .B2(new_n498), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n500), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n493), .A2(new_n498), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n510), .A3(new_n509), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n480), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n516), .A4(new_n518), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n511), .A2(new_n499), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n518), .B(KEYINPUT13), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n520), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT11), .B(G169gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n528), .B(new_n529), .Z(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n531), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n520), .A2(new_n533), .A3(new_n521), .A4(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n479), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT92), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(new_n548), .A3(G85gat), .A4(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(G99gat), .ZN(new_n550));
  INV_X1    g349(.A(G106gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT8), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G99gat), .B(G106gat), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(new_n549), .A3(new_n552), .A4(new_n545), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n500), .A2(new_n513), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n557), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n515), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n540), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(new_n562), .A3(new_n540), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n567), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G71gat), .B(G78gat), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G64gat), .ZN(new_n579));
  INV_X1    g378(.A(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G57gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT88), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n581), .A3(KEYINPUT88), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n576), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n579), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n581), .B(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n577), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT21), .ZN(new_n593));
  AND2_X1   g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G127gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n591), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n584), .A2(new_n585), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n576), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT91), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n511), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n596), .A2(new_n604), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n347), .ZN(new_n610));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n574), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n555), .A2(new_n618), .A3(new_n557), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n599), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n558), .ZN(new_n621));
  AOI21_X1  g420(.A(KEYINPUT10), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n558), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n600), .A2(new_n602), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G230gat), .ZN(new_n626));
  OAI22_X1  g425(.A1(new_n622), .A2(new_n625), .B1(new_n626), .B2(new_n271), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n271), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n620), .A2(new_n628), .A3(new_n621), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT96), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n616), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n536), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n405), .A2(new_n410), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n411), .B1(new_n645), .B2(new_n404), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n476), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(KEYINPUT42), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n652), .B(new_n653), .C1(new_n508), .C2(new_n649), .ZN(G1325gat));
  AND3_X1   g453(.A1(new_n295), .A2(KEYINPUT36), .A3(new_n299), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT36), .B1(new_n295), .B2(new_n299), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n644), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n295), .A2(new_n299), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(G15gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n644), .B2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n644), .A2(new_n466), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n614), .A2(new_n615), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n574), .A3(new_n642), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT98), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n536), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n646), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n483), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(new_n535), .ZN(new_n674));
  INV_X1    g473(.A(new_n642), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n666), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT99), .B1(new_n466), .B2(new_n469), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n646), .A2(new_n476), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT81), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n437), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n432), .A2(new_n436), .A3(KEYINPUT81), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n463), .A2(new_n685), .B1(new_n474), .B2(new_n478), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n686), .A2(new_n574), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(new_n479), .B2(new_n574), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n676), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n646), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n692), .ZN(G1328gat));
  NOR2_X1   g492(.A1(new_n476), .A2(new_n490), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n670), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  OAI21_X1  g495(.A(new_n490), .B1(new_n691), .B2(new_n476), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n691), .B2(new_n657), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT47), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n670), .A2(new_n702), .A3(new_n659), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n701), .B(new_n704), .ZN(G1330gat));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n670), .A2(new_n706), .A3(new_n682), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  OAI21_X1  g507(.A(G50gat), .B1(new_n691), .B2(new_n437), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(KEYINPUT102), .B2(KEYINPUT48), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n706), .A2(KEYINPUT48), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n691), .B2(new_n466), .ZN(new_n713));
  AOI22_X1  g512(.A1(KEYINPUT48), .A2(new_n710), .B1(new_n711), .B2(new_n713), .ZN(G1331gat));
  NAND3_X1  g513(.A1(new_n616), .A2(new_n674), .A3(new_n675), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n454), .A2(new_n458), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n454), .A2(new_n446), .A3(new_n458), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n406), .A2(new_n408), .B1(new_n441), .B2(new_n443), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n472), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n439), .A2(new_n403), .A3(new_n402), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n411), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(new_n343), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n657), .A2(new_n724), .A3(new_n677), .A4(new_n684), .ZN(new_n725));
  OAI21_X1  g524(.A(KEYINPUT35), .B1(new_n475), .B2(new_n678), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n473), .A2(new_n723), .A3(new_n471), .A4(new_n476), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n715), .B1(new_n725), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n671), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n444), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT49), .B(G64gat), .Z(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g534(.A(new_n657), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(G71gat), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT103), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n729), .A2(new_n659), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(G71gat), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n729), .A2(new_n682), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n666), .A2(new_n535), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n675), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n479), .A2(new_n574), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n573), .B1(new_n725), .B2(new_n728), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n687), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n671), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G85gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n686), .A2(new_n574), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n574), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(KEYINPUT51), .A3(new_n744), .A4(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n744), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n753), .B2(new_n754), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(KEYINPUT105), .A3(KEYINPUT51), .A4(new_n756), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n744), .B1(new_n748), .B2(KEYINPUT104), .ZN(new_n764));
  INV_X1    g563(.A(new_n756), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n759), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n675), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n646), .A2(G85gat), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n752), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NOR2_X1   g569(.A1(new_n476), .A2(G92gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n675), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(G92gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n750), .B2(new_n444), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n675), .A2(new_n771), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n766), .B2(new_n757), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT106), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(KEYINPUT52), .C1(new_n778), .C2(new_n774), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n780), .A3(new_n782), .ZN(G1337gat));
  NAND2_X1  g582(.A1(new_n750), .A2(new_n736), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n550), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n785), .B2(new_n784), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n659), .A2(new_n550), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n768), .B2(new_n788), .ZN(G1338gat));
  INV_X1    g588(.A(new_n745), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n682), .B(new_n790), .C1(new_n688), .C2(new_n690), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G106gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(KEYINPUT108), .A3(G106gat), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n766), .A2(new_n757), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n642), .A2(G106gat), .A3(new_n437), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT109), .Z(new_n798));
  OAI211_X1 g597(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n767), .A2(new_n797), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n472), .B(new_n790), .C1(new_n688), .C2(new_n690), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n551), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n750), .A2(KEYINPUT110), .A3(new_n472), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT53), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n800), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n620), .A2(new_n621), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n623), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n600), .A2(new_n602), .A3(new_n624), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n628), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n814), .A2(new_n627), .A3(KEYINPUT54), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n634), .B1(new_n627), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n810), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n628), .B1(new_n812), .B2(new_n813), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n636), .B1(new_n820), .B2(new_n816), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n627), .A3(KEYINPUT54), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n637), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n523), .A2(new_n524), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n517), .A2(new_n519), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n517), .A2(KEYINPUT112), .A3(new_n519), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n530), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n574), .A3(new_n534), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n809), .B1(new_n824), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n823), .A2(new_n637), .ZN(new_n834));
  INV_X1    g633(.A(new_n530), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n828), .B2(new_n829), .ZN(new_n836));
  INV_X1    g635(.A(new_n534), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n836), .A2(new_n837), .A3(new_n573), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n834), .A2(new_n838), .A3(KEYINPUT113), .A4(new_n819), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n836), .A2(new_n837), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n640), .A2(new_n841), .A3(new_n641), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n819), .A2(new_n535), .A3(new_n637), .A4(new_n823), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n574), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n667), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n616), .A2(new_n674), .A3(new_n642), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n682), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n646), .A2(new_n444), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n660), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851), .B2(new_n674), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n646), .B1(new_n845), .B2(new_n846), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n475), .A2(new_n444), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n535), .A2(new_n255), .A3(new_n256), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(G1340gat));
  OR3_X1    g656(.A1(new_n855), .A2(G120gat), .A3(new_n642), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n847), .A2(new_n675), .A3(new_n850), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G120gat), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(KEYINPUT114), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT115), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n851), .B2(new_n667), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n666), .A2(new_n248), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n855), .B2(new_n866), .ZN(G1342gat));
  NAND4_X1  g666(.A1(new_n853), .A2(new_n246), .A3(new_n574), .A4(new_n854), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n851), .B2(new_n573), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n736), .A2(new_n849), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n437), .B1(new_n845), .B2(new_n846), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n682), .A2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n823), .A2(new_n637), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT55), .B1(new_n821), .B2(new_n822), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n819), .A2(KEYINPUT117), .A3(new_n637), .A4(new_n823), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n535), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n574), .B1(new_n885), .B2(new_n842), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n667), .B1(new_n886), .B2(new_n840), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n879), .B1(new_n887), .B2(new_n846), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n535), .B(new_n874), .C1(new_n878), .C2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT58), .B1(new_n889), .B2(G141gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n736), .A2(new_n437), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n845), .A2(new_n846), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n671), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n674), .A2(G141gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n853), .A2(KEYINPUT118), .A3(new_n891), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n895), .A2(new_n476), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n444), .B1(new_n893), .B2(new_n894), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n896), .A4(new_n897), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n890), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n889), .A2(G141gat), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n853), .A2(new_n476), .A3(new_n891), .A4(new_n896), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n873), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n907), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n899), .A3(new_n902), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n911), .ZN(G1344gat));
  AND2_X1   g711(.A1(new_n900), .A2(new_n897), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n675), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n674), .B1(new_n824), .B2(new_n880), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n917), .A2(new_n884), .B1(new_n675), .B2(new_n841), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n918), .A2(new_n574), .B1(new_n824), .B2(new_n832), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n919), .A2(new_n667), .B1(new_n674), .B2(new_n643), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n466), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n824), .A2(new_n832), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n667), .B1(new_n886), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n846), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT121), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n875), .A2(new_n877), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n675), .B(new_n874), .C1(new_n927), .C2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n916), .B1(new_n930), .B2(G148gat), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n878), .A2(new_n888), .ZN(new_n932));
  INV_X1    g731(.A(new_n874), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI211_X1 g733(.A(KEYINPUT59), .B(new_n914), .C1(new_n934), .C2(new_n675), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n915), .B1(new_n931), .B2(new_n935), .ZN(G1345gat));
  AOI21_X1  g735(.A(G155gat), .B1(new_n913), .B2(new_n666), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n666), .A2(G155gat), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n934), .B2(new_n939), .ZN(G1346gat));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n574), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n348), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n913), .A2(new_n348), .A3(new_n574), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1347gat));
  NAND2_X1  g745(.A1(new_n646), .A2(new_n444), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n660), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n847), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G169gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n950), .A2(new_n951), .A3(new_n674), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n671), .B1(new_n845), .B2(new_n846), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n475), .A2(new_n476), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n535), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n952), .B1(new_n951), .B2(new_n957), .ZN(G1348gat));
  OAI21_X1  g757(.A(G176gat), .B1(new_n950), .B2(new_n642), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n642), .A2(G176gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n955), .B2(new_n960), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n950), .B2(new_n667), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n666), .A2(new_n217), .A3(new_n218), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n955), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n964), .B(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n956), .A2(new_n219), .A3(new_n574), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n847), .A2(new_n574), .A3(new_n949), .ZN(new_n968));
  XNOR2_X1  g767(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n968), .A2(G190gat), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n968), .B2(G190gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1351gat));
  AND3_X1   g771(.A1(new_n953), .A2(new_n444), .A3(new_n891), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n535), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n736), .A2(new_n948), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n922), .A2(new_n926), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT57), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n976), .B1(new_n979), .B2(new_n928), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n535), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  INV_X1    g781(.A(G204gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n973), .A2(new_n983), .A3(new_n675), .ZN(new_n984));
  XOR2_X1   g783(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n985));
  XNOR2_X1  g784(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AOI211_X1 g785(.A(new_n642), .B(new_n976), .C1(new_n979), .C2(new_n928), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n983), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n317), .A3(new_n666), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n666), .B(new_n975), .C1(new_n927), .C2(new_n929), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n318), .A3(new_n574), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n980), .A2(new_n574), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(new_n318), .ZN(G1355gat));
endmodule


