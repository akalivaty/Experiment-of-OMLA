//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n475), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(new_n471), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n465), .A2(new_n474), .A3(new_n479), .ZN(G160));
  OAI21_X1  g055(.A(KEYINPUT69), .B1(new_n470), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n458), .A2(new_n482), .A3(new_n460), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n464), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(KEYINPUT70), .A2(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT70), .A2(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n460), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n493), .A2(new_n494), .B1(new_n470), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n464), .A2(new_n458), .A3(G138), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n458), .A3(new_n499), .A4(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OR3_X1    g083(.A1(new_n507), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n510), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(G543), .ZN(new_n516));
  AND3_X1   g091(.A1(new_n506), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n507), .B2(new_n508), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n509), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT73), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n502), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n525), .ZN(G166));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n517), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n527), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(new_n517), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n521), .A2(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n546), .A2(G651), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n517), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT75), .Z(G188));
  NAND3_X1  g133(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n517), .A2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n502), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G166), .ZN(G303));
  OAI21_X1  g143(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n517), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n527), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n517), .A2(G86), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n503), .A2(new_n505), .A3(G48), .A4(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT76), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n515), .A2(G61), .A3(new_n516), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n502), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n502), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n527), .A2(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n539), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n527), .A2(G54), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n502), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n517), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G321));
  NOR2_X1   g173(.A1(new_n565), .A2(G868), .ZN(new_n599));
  AND2_X1   g174(.A1(G286), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT78), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(KEYINPUT78), .B2(new_n600), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(KEYINPUT78), .B2(new_n600), .ZN(G280));
  XOR2_X1   g178(.A(KEYINPUT79), .B(G559), .Z(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(G860), .B2(new_n604), .ZN(G148));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n604), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT80), .Z(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n458), .A2(new_n473), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2100), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n486), .A2(G123), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n484), .A2(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n615), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(KEYINPUT14), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT83), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n632), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2072), .B(G2078), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n642), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n647), .A2(KEYINPUT17), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n647), .B2(KEYINPUT17), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n648), .A2(new_n649), .A3(new_n643), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  OAI221_X1 g238(.A(new_n659), .B1(new_n656), .B2(new_n660), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1991), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OR3_X1    g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(G229));
  INV_X1    g250(.A(G29), .ZN(new_n676));
  NOR2_X1   g251(.A1(G162), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(G35), .ZN(new_n678));
  OAI21_X1  g253(.A(KEYINPUT102), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(KEYINPUT102), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G2090), .Z(new_n683));
  INV_X1    g258(.A(G19), .ZN(new_n684));
  OAI21_X1  g259(.A(KEYINPUT88), .B1(new_n684), .B2(G16), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n684), .A2(KEYINPUT88), .A3(G16), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n686), .C1(new_n551), .C2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(G1341), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n484), .A2(G141), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT97), .ZN(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT98), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n486), .A2(G129), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n473), .A2(G105), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n693), .A2(KEYINPUT26), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT99), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(new_n676), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n676), .B2(G32), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n683), .A2(new_n689), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n676), .A2(G26), .ZN(new_n708));
  INV_X1    g283(.A(new_n486), .ZN(new_n709));
  INV_X1    g284(.A(G128), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n709), .A2(KEYINPUT89), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT89), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n466), .B1(new_n713), .B2(KEYINPUT90), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n714), .B1(KEYINPUT90), .B2(new_n713), .C1(G116), .C2(new_n464), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n711), .B(new_n716), .C1(G140), .C2(new_n484), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(new_n676), .ZN(new_n718));
  MUX2_X1   g293(.A(new_n708), .B(new_n718), .S(KEYINPUT28), .Z(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(G2067), .ZN(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G171), .B2(G16), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(G1961), .ZN(new_n723));
  NOR2_X1   g298(.A1(G29), .A2(G33), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT91), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT92), .B(KEYINPUT93), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT25), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n484), .A2(G139), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n464), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n727), .A2(new_n728), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(new_n676), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n676), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n676), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AND4_X1   g316(.A1(new_n720), .A2(new_n723), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n687), .A2(G20), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT23), .B1(new_n565), .B2(new_n687), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n743), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n676), .B1(new_n750), .B2(G34), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(new_n750), .B2(G34), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n752), .B2(new_n751), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT96), .Z(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n719), .A2(G2067), .B1(G2084), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n735), .A2(new_n736), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n756), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n742), .A2(new_n748), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G286), .A2(new_n687), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT100), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G16), .B2(G21), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n722), .A2(G1961), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT31), .B(G11), .Z(new_n771));
  XOR2_X1   g346(.A(KEYINPUT101), .B(KEYINPUT30), .Z(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(G28), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n770), .B(new_n775), .C1(new_n676), .C2(new_n620), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n768), .A2(new_n769), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n596), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n781), .C1(new_n705), .C2(new_n704), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n707), .A2(new_n763), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n687), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n687), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1971), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n687), .A2(G6), .ZN(new_n787));
  INV_X1    g362(.A(G305), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n687), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G23), .B(G288), .S(G16), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT86), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n786), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n587), .A2(new_n687), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n687), .B2(G24), .ZN(new_n802));
  INV_X1    g377(.A(G1986), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n676), .A2(G25), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n807));
  INV_X1    g382(.A(G119), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n709), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G131), .B2(new_n484), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n806), .B1(new_n810), .B2(new_n676), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  NOR3_X1   g388(.A1(new_n804), .A2(new_n805), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n799), .A2(new_n800), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(KEYINPUT87), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n783), .A2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  INV_X1    g395(.A(G860), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n596), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n517), .A2(G93), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n502), .ZN(new_n827));
  AOI211_X1 g402(.A(new_n825), .B(new_n827), .C1(G55), .C2(new_n527), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n550), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n824), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT105), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n821), .B1(KEYINPUT39), .B2(new_n831), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n828), .A2(new_n821), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n620), .B(G162), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G160), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT112), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n484), .A2(G142), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT108), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n464), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n845), .A2(new_n847), .B1(new_n486), .B2(G130), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n810), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT109), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n613), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT111), .ZN(new_n853));
  MUX2_X1   g428(.A(new_n702), .B(new_n700), .S(new_n734), .Z(new_n854));
  AOI211_X1 g429(.A(KEYINPUT107), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n498), .A2(new_n500), .ZN(new_n857));
  INV_X1    g432(.A(new_n496), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n717), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n842), .B1(new_n853), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n852), .A2(new_n862), .A3(KEYINPUT111), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT110), .B(G37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n852), .ZN(new_n868));
  INV_X1    g443(.A(new_n613), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n851), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n862), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n841), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n867), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT40), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n866), .A2(new_n875), .A3(new_n867), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G395));
  NAND2_X1  g452(.A1(new_n608), .A2(new_n830), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n607), .A2(new_n829), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n596), .A2(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n593), .A2(new_n595), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n565), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n881), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n881), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n878), .B(new_n879), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n587), .B(G288), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G303), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n788), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n884), .A2(new_n889), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n884), .B2(new_n889), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G868), .B2(new_n828), .ZN(G295));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n828), .ZN(G331));
  XOR2_X1   g473(.A(G286), .B(G171), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n829), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n881), .B2(new_n883), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n886), .A2(new_n888), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n901), .B(new_n892), .C1(new_n902), .C2(new_n900), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n867), .A3(new_n907), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT44), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n908), .A2(new_n909), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n909), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  OAI211_X1 g494(.A(KEYINPUT45), .B(new_n919), .C1(new_n855), .C2(new_n859), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n465), .A2(new_n474), .A3(G40), .A4(new_n479), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n857), .A2(new_n858), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT56), .B(G2072), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT57), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n562), .B2(new_n564), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n563), .A2(new_n502), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(KEYINPUT57), .A3(new_n561), .A4(new_n560), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n922), .A2(new_n933), .A3(new_n919), .ZN(new_n934));
  INV_X1    g509(.A(new_n921), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(KEYINPUT118), .B(G1956), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT119), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT119), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n927), .A2(new_n932), .A3(new_n939), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT121), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT61), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT61), .B1(new_n941), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n927), .A2(new_n939), .ZN(new_n949));
  INV_X1    g524(.A(new_n932), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT121), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT120), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n937), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(KEYINPUT120), .ZN(new_n956));
  AOI21_X1  g531(.A(G1348), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(G164), .A2(G1384), .ZN(new_n959));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n935), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(KEYINPUT60), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT60), .ZN(new_n963));
  INV_X1    g538(.A(new_n961), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n596), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n920), .A2(new_n925), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT58), .B(G1341), .Z(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n923), .B2(new_n921), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n550), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT59), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n958), .A2(KEYINPUT60), .A3(new_n882), .A4(new_n961), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n966), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n882), .B1(new_n958), .B2(new_n961), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n950), .B2(new_n949), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n953), .A2(new_n975), .B1(new_n977), .B2(new_n944), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n922), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n924), .B1(G164), .B2(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n935), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n767), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n761), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT122), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT51), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n937), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n988), .A2(new_n761), .B1(new_n982), .B2(new_n767), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n979), .B1(new_n989), .B2(G168), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n985), .ZN(new_n992));
  NAND2_X1  g567(.A1(G286), .A2(G8), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n986), .A3(KEYINPUT51), .A4(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n989), .A2(new_n993), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(KEYINPUT116), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(G166), .B2(new_n979), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT55), .B(G8), .C1(new_n520), .C2(new_n525), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n935), .A2(new_n981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G164), .A2(new_n856), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n1006), .A2(G1971), .B1(G2090), .B2(new_n937), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1001), .B1(new_n1007), .B2(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1971), .B1(new_n920), .B2(new_n925), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n937), .A2(G2090), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1001), .B(G8), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n997), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n955), .A2(new_n956), .ZN(new_n1014));
  INV_X1    g589(.A(G1961), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n920), .A2(new_n925), .A3(new_n740), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n925), .A2(KEYINPUT53), .A3(new_n740), .A4(new_n980), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n1022));
  XNOR2_X1  g597(.A(G171), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n919), .B1(new_n855), .B2(new_n859), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT45), .B1(new_n1024), .B2(KEYINPUT113), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1005), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n740), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT123), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n471), .B1(new_n459), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n477), .A2(KEYINPUT123), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n474), .B(new_n1029), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1023), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1014), .A2(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1021), .A2(new_n1023), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n576), .B2(new_n580), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n573), .A2(new_n575), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1041), .A2(G1981), .A3(new_n579), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n979), .B1(new_n935), .B2(new_n959), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n576), .A2(new_n1039), .A3(new_n580), .ZN(new_n1045));
  OAI21_X1  g620(.A(G1981), .B1(new_n1041), .B2(new_n579), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT49), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1044), .ZN(new_n1049));
  INV_X1    g624(.A(G1976), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G288), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT52), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1050), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1044), .B(new_n1053), .C1(new_n1050), .C2(G288), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1048), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT116), .B(G8), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n996), .A2(new_n1013), .A3(new_n1037), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n997), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1001), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1064), .B2(new_n1011), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT124), .A3(new_n996), .A4(new_n1037), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n978), .A2(new_n1060), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n985), .A2(G168), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1072), .B2(KEYINPUT63), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1071), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1013), .A2(new_n1057), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1075), .A2(KEYINPUT117), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT63), .A3(new_n1055), .A4(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(G1976), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1049), .B1(new_n1083), .B2(new_n1045), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1012), .B2(new_n1055), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT115), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1069), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1069), .A2(new_n1080), .A3(new_n1086), .A4(KEYINPUT125), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n1092));
  AOI21_X1  g667(.A(G301), .B1(new_n1036), .B2(new_n1020), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(new_n1067), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1028), .A2(new_n921), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G290), .A2(G1986), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n587), .A2(new_n803), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1096), .B(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n717), .B(new_n960), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1096), .A2(new_n967), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1101), .A2(new_n1102), .B1(new_n702), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n810), .B(new_n812), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1101), .A2(G1996), .A3(new_n700), .ZN(new_n1108));
  AND4_X1   g683(.A1(new_n1099), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1095), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT48), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1103), .B(KEYINPUT46), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n700), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1117), .A2(KEYINPUT47), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(KEYINPUT47), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n810), .A2(new_n812), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT126), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1105), .A2(new_n1108), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n717), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(G2067), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1101), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1110), .A2(new_n1126), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g702(.A(G319), .ZN(new_n1129));
  NOR3_X1   g703(.A1(G401), .A2(new_n1129), .A3(G227), .ZN(new_n1130));
  NAND4_X1  g704(.A1(new_n673), .A2(KEYINPUT127), .A3(new_n674), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n673), .A2(new_n674), .A3(new_n1130), .ZN(new_n1132));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n1133));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g708(.A1(new_n864), .A2(new_n865), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n872), .A2(new_n867), .ZN(new_n1136));
  OAI211_X1 g710(.A(new_n1131), .B(new_n1134), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n914), .A2(new_n916), .ZN(new_n1138));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n1138), .ZN(G308));
  AND2_X1   g713(.A1(new_n1134), .A2(new_n1131), .ZN(new_n1140));
  NAND4_X1  g714(.A1(new_n1140), .A2(new_n873), .A3(new_n916), .A4(new_n914), .ZN(G225));
endmodule


