//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT68), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT69), .Z(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n469), .A2(G137), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n475));
  OAI211_X1 g050(.A(G101), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(KEYINPUT71), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT71), .B1(new_n473), .B2(new_n476), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n480), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n470), .ZN(new_n482));
  NOR3_X1   g057(.A1(new_n478), .A2(new_n479), .A3(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n469), .A2(new_n472), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT73), .Z(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n469), .A2(G126), .A3(new_n472), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n470), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n470), .A2(G138), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT4), .B1(new_n480), .B2(new_n502), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT74), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(G88), .B1(new_n513), .B2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n509), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT75), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(G166));
  XOR2_X1   g099(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT76), .B(G51), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n513), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n510), .A2(G543), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT78), .B(G52), .Z(new_n539));
  OAI22_X1  g114(.A1(new_n511), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n512), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n535), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n513), .A2(G53), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n535), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n512), .A2(G91), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(G166), .ZN(G303));
  INV_X1    g133(.A(G87), .ZN(new_n559));
  INV_X1    g134(.A(G49), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n511), .A2(new_n559), .B1(new_n538), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G288));
  NAND3_X1  g140(.A1(new_n509), .A2(G86), .A3(new_n510), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n508), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT5), .B1(KEYINPUT74), .B2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(G61), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n535), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(G72), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G60), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n516), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n535), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n579), .B2(new_n578), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n512), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n512), .A2(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n516), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n584), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G299), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G297));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g179(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n605));
  INV_X1    g180(.A(new_n480), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n487), .A2(G123), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n612), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G135), .B2(new_n485), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n610), .A2(new_n616), .ZN(G156));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2438), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2430), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n621), .B2(new_n620), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n623), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(G14), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT80), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT18), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(KEYINPUT17), .ZN(new_n640));
  INV_X1    g215(.A(new_n634), .ZN(new_n641));
  INV_X1    g216(.A(new_n635), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n641), .A2(new_n637), .A3(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT82), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT81), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n651));
  XNOR2_X1  g226(.A(G1971), .B(G1976), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n656), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n658), .B(new_n661), .C1(new_n653), .C2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(G229));
  XNOR2_X1  g246(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT95), .ZN(new_n673));
  NAND3_X1  g248(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OAI211_X1 g250(.A(G105), .B(new_n470), .C1(new_n474), .C2(new_n475), .ZN(new_n676));
  AOI22_X1  g251(.A1(G129), .A2(new_n487), .B1(new_n485), .B2(G141), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(G32), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT27), .B(G1996), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n485), .A2(G139), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT25), .Z(new_n686));
  AOI22_X1  g261(.A1(new_n480), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n684), .B(new_n686), .C1(new_n470), .C2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(G33), .B(new_n688), .S(G29), .Z(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2072), .Z(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(G168), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(G21), .ZN(new_n693));
  INV_X1    g268(.A(G1966), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT31), .B(G11), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT30), .B(G28), .Z(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G29), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n693), .B2(new_n694), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n683), .A2(new_n690), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G19), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n701), .A2(KEYINPUT89), .A3(G16), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT89), .B1(new_n701), .B2(G16), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n702), .B(new_n703), .C1(new_n545), .C2(new_n691), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1341), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n679), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  OR2_X1    g282(.A1(G104), .A2(G2105), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n708), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT90), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G140), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n487), .A2(G128), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n707), .B1(new_n714), .B2(new_n679), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT91), .B(G2067), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n615), .A2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n705), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n691), .A2(G5), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G171), .B2(new_n691), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1961), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n691), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT102), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT23), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G299), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1956), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR4_X1   g305(.A1(new_n700), .A2(new_n720), .A3(new_n724), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n494), .A2(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n679), .A2(G35), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT99), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n735));
  AND3_X1   g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n732), .B2(new_n734), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n736), .A2(new_n737), .A3(G2090), .ZN(new_n738));
  NOR2_X1   g313(.A1(G4), .A2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT88), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n587), .A2(new_n591), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n691), .ZN(new_n742));
  INV_X1    g317(.A(G1348), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G27), .A2(G29), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G164), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2078), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n731), .A2(new_n738), .A3(new_n748), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n681), .A2(new_n682), .B1(G1961), .B2(new_n722), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G160), .B2(new_n679), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT92), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G2084), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(G2084), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(G2090), .B1(new_n736), .B2(new_n737), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT101), .Z(new_n765));
  NOR3_X1   g340(.A1(new_n749), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G166), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G16), .B2(G22), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT86), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(KEYINPUT86), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G1971), .ZN(new_n772));
  INV_X1    g347(.A(G1971), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n769), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G23), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n512), .A2(G87), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n513), .A2(G49), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n776), .A2(KEYINPUT85), .A3(new_n777), .A4(new_n562), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n561), .B2(new_n563), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n782), .B(new_n783), .Z(new_n784));
  NOR2_X1   g359(.A1(G6), .A2(G16), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n574), .B2(G16), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1981), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n772), .A2(new_n774), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  MUX2_X1   g366(.A(G24), .B(G290), .S(G16), .Z(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G1986), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n487), .A2(G119), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT84), .B1(G95), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(KEYINPUT84), .A2(G95), .A3(G2105), .ZN(new_n798));
  OAI221_X1 g373(.A(G2104), .B1(G107), .B2(new_n470), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G25), .B(new_n800), .S(G29), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT35), .B(G1991), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n792), .A2(G1986), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n793), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n790), .B2(KEYINPUT34), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n791), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n791), .B2(new_n806), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n766), .B1(new_n808), .B2(new_n809), .ZN(G150));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n811));
  XNOR2_X1  g386(.A(G150), .B(new_n811), .ZN(G311));
  NAND2_X1  g387(.A1(new_n592), .A2(G559), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT38), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT104), .B(G93), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n511), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(new_n535), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n816), .B(new_n818), .C1(G55), .C2(new_n513), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n545), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n814), .B(new_n820), .Z(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n819), .A2(new_n823), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  XOR2_X1   g403(.A(KEYINPUT107), .B(G37), .Z(new_n829));
  INV_X1    g404(.A(KEYINPUT106), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n688), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT105), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G164), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n487), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n470), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G142), .B2(new_n485), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n608), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n678), .B(new_n714), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n800), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n615), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G162), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n842), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n843), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n843), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n829), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g426(.A(new_n820), .B(new_n601), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n592), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n596), .A2(new_n741), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n858));
  OR3_X1    g433(.A1(new_n855), .A2(KEYINPUT109), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT109), .B1(new_n855), .B2(new_n858), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n853), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n596), .A2(new_n741), .A3(KEYINPUT108), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n859), .B(new_n860), .C1(new_n864), .C2(KEYINPUT41), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n852), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT110), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(KEYINPUT110), .A3(new_n852), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT42), .ZN(new_n871));
  XNOR2_X1  g446(.A(G166), .B(G290), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n781), .B(G305), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n875), .A3(new_n869), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  OAI21_X1  g453(.A(G868), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n819), .A2(G868), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(G295));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT111), .ZN(new_n883));
  AOI21_X1  g458(.A(G286), .B1(new_n883), .B2(G171), .ZN(new_n884));
  NAND2_X1  g459(.A1(G301), .A2(KEYINPUT111), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n820), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n820), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n855), .A2(new_n858), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT113), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n864), .A2(KEYINPUT41), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT114), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n887), .A2(KEYINPUT112), .A3(new_n888), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n886), .A2(new_n820), .A3(KEYINPUT112), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n856), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n874), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n896), .A2(new_n897), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n901), .A2(new_n865), .B1(new_n855), .B2(new_n889), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n874), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n829), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n900), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n902), .A2(new_n874), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n902), .B2(new_n874), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT43), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT43), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(new_n914), .ZN(G397));
  XNOR2_X1  g490(.A(new_n678), .B(G1996), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n713), .B(G2067), .Z(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n800), .B(new_n802), .Z(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(G164), .B2(G1384), .ZN(new_n922));
  INV_X1    g497(.A(new_n479), .ZN(new_n923));
  INV_X1    g498(.A(new_n482), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(G40), .A3(new_n924), .A4(new_n477), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n927), .A2(G1986), .A3(G290), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n794), .A2(new_n795), .A3(new_n802), .A4(new_n799), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n918), .A2(new_n933), .B1(G2067), .B2(new_n713), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n926), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n927), .B1(new_n917), .B2(new_n678), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n932), .B(new_n935), .C1(new_n936), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n936), .B2(new_n942), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n778), .A2(new_n780), .A3(G1976), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  INV_X1    g521(.A(new_n503), .ZN(new_n947));
  INV_X1    g522(.A(new_n500), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT70), .B(G2104), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n471), .B1(new_n949), .B2(KEYINPUT3), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n948), .B1(new_n950), .B2(G126), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n951), .B2(new_n470), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n946), .B1(new_n952), .B2(new_n498), .ZN(new_n953));
  OAI211_X1 g528(.A(G8), .B(new_n945), .C1(new_n953), .C2(new_n925), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n954), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n564), .B2(G1976), .ZN(new_n957));
  OAI21_X1  g532(.A(G8), .B1(new_n953), .B2(new_n925), .ZN(new_n958));
  OAI21_X1  g533(.A(G1981), .B1(new_n568), .B2(new_n573), .ZN(new_n959));
  INV_X1    g534(.A(G61), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n507), .B2(new_n508), .ZN(new_n961));
  INV_X1    g536(.A(new_n572), .ZN(new_n962));
  OAI21_X1  g537(.A(G651), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1981), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n566), .A4(new_n567), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n965), .A3(KEYINPUT49), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI22_X1  g545(.A1(new_n954), .A2(new_n957), .B1(new_n958), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT115), .B1(new_n954), .B2(KEYINPUT52), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n955), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  INV_X1    g549(.A(G40), .ZN(new_n975));
  NOR4_X1   g550(.A1(new_n478), .A2(new_n479), .A3(new_n975), .A4(new_n482), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n499), .A2(new_n500), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n503), .B1(new_n977), .B2(G2105), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n496), .A2(new_n497), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n470), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n922), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n694), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n986), .A3(new_n946), .ZN(new_n987));
  INV_X1    g562(.A(G2084), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n976), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n974), .B(G286), .C1(new_n984), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n773), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n925), .B1(new_n953), .B2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(G2090), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n521), .A2(new_n523), .A3(G8), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(G8), .A3(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n973), .A2(new_n990), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n974), .B1(new_n991), .B2(new_n994), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n998), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n996), .B(KEYINPUT55), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n985), .A2(new_n976), .A3(new_n987), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n1005), .A2(new_n993), .B1(new_n983), .B2(new_n773), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT116), .B(new_n1004), .C1(new_n1006), .C2(new_n974), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1000), .A2(KEYINPUT117), .A3(new_n1003), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT63), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n973), .A2(new_n990), .A3(new_n999), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1008), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1000), .B(KEYINPUT63), .C1(new_n998), .C2(new_n1002), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(G1976), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n958), .B2(new_n970), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n958), .B1(new_n1018), .B2(new_n965), .ZN(new_n1019));
  INV_X1    g594(.A(new_n999), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n973), .ZN(new_n1021));
  OR4_X1    g596(.A1(KEYINPUT118), .A2(new_n953), .A3(new_n925), .A4(G2067), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n985), .A2(new_n976), .A3(new_n987), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n743), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n978), .B2(new_n980), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n976), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n1026), .B2(G2067), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n976), .B1(new_n986), .B2(new_n1025), .ZN(new_n1029));
  NOR3_X1   g604(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n729), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G299), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n552), .A2(KEYINPUT57), .A3(new_n554), .A4(new_n555), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT56), .B(G2072), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n922), .A2(new_n982), .A3(new_n976), .A4(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1028), .A2(new_n1038), .A3(new_n592), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1035), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1956), .B1(new_n992), .B2(new_n987), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1037), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT60), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1028), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1022), .A2(new_n1024), .A3(KEYINPUT60), .A4(new_n1027), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n592), .A3(new_n1047), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n1028), .A2(new_n1045), .A3(new_n592), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1031), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1035), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1051), .A2(new_n1052), .A3(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1043), .B2(new_n1038), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT58), .B(G1341), .Z(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n953), .B2(new_n925), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT119), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1026), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n922), .A2(new_n982), .A3(new_n939), .A4(new_n976), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1056), .B1(new_n1063), .B2(new_n545), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(new_n1056), .A3(new_n545), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1053), .A2(new_n1055), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1066), .B2(KEYINPUT120), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  OAI221_X1 g643(.A(new_n1068), .B1(new_n1064), .B2(new_n1065), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1044), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n983), .B2(G2078), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1023), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1071), .A2(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n922), .A2(new_n982), .A3(new_n976), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n481), .A2(KEYINPUT125), .ZN(new_n1082));
  OAI21_X1  g657(.A(G2105), .B1(new_n481), .B2(KEYINPUT125), .ZN(new_n1083));
  OAI211_X1 g658(.A(G40), .B(new_n1075), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n478), .A2(new_n479), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(KEYINPUT124), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1085), .A2(KEYINPUT124), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n922), .A4(new_n982), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1072), .A2(new_n1074), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1080), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1003), .A2(new_n1007), .A3(new_n999), .A4(new_n973), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(G171), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1072), .A2(G301), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1095), .A2(KEYINPUT54), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n984), .A2(G168), .A3(new_n989), .ZN(new_n1099));
  AND2_X1   g674(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1103), .A3(new_n1100), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n974), .B1(new_n984), .B2(new_n989), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G286), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT122), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1101), .A2(KEYINPUT51), .B1(G286), .B2(new_n1105), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1104), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1093), .B(new_n1098), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1016), .B(new_n1021), .C1(new_n1070), .C2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT62), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1107), .A2(KEYINPUT122), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n1109), .A3(new_n1104), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1094), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT126), .A3(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n1108), .C2(new_n1111), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1116), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1113), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(G290), .B(G1986), .Z(new_n1129));
  AOI21_X1  g704(.A(new_n927), .B1(new_n920), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n944), .B1(new_n1128), .B2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g706(.A1(G401), .A2(new_n463), .A3(G227), .ZN(new_n1133));
  OAI21_X1  g707(.A(new_n1133), .B1(new_n669), .B2(new_n670), .ZN(new_n1134));
  INV_X1    g708(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g709(.A(new_n850), .B(new_n1135), .C1(new_n912), .C2(new_n913), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


