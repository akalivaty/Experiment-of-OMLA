//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT81), .A2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(G237), .A2(G953), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(G214), .C1(KEYINPUT81), .C2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n197), .A3(KEYINPUT82), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT18), .A2(G131), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT72), .A2(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT72), .A2(G125), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(G125), .A2(G140), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  XOR2_X1   g021(.A(G125), .B(G140), .Z(new_n208));
  OR2_X1    g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n195), .A2(new_n197), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(G131), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n213), .A2(KEYINPUT17), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT72), .A2(G125), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT72), .A2(G125), .ZN(new_n218));
  OAI21_X1  g032(.A(G140), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n205), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n201), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n202), .B2(new_n203), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n215), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT16), .B1(new_n204), .B2(new_n205), .ZN(new_n225));
  INV_X1    g039(.A(new_n223), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(G146), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n228));
  AND4_X1   g042(.A1(new_n228), .A2(new_n212), .A3(KEYINPUT17), .A4(G131), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n195), .B2(new_n197), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n231), .B2(KEYINPUT17), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n224), .B(new_n227), .C1(new_n229), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n214), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(G146), .B1(new_n225), .B2(new_n226), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n221), .A2(new_n215), .A3(new_n223), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT84), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n231), .A2(new_n228), .A3(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT85), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n190), .B(new_n211), .C1(new_n235), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(new_n234), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT85), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n214), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n190), .B1(new_n248), .B2(new_n211), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n187), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G475), .ZN(new_n251));
  INV_X1    g065(.A(G478), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT15), .ZN(new_n253));
  XNOR2_X1  g067(.A(G128), .B(G143), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G116), .B(G122), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT14), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G116), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT14), .A3(G122), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(G107), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G107), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT87), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT87), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n257), .A2(new_n266), .A3(new_n263), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n256), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G128), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n270), .B(G134), .C1(new_n272), .C2(new_n269), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n257), .B(new_n263), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n255), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT9), .B(G234), .ZN(new_n278));
  INV_X1    g092(.A(G217), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n278), .A2(new_n279), .A3(G953), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n268), .A2(new_n276), .A3(new_n280), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT70), .B(G902), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT88), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n268), .A2(new_n276), .A3(new_n280), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n280), .B1(new_n268), .B2(new_n276), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT88), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n253), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n285), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n282), .B2(new_n283), .ZN(new_n293));
  OAI22_X1  g107(.A1(new_n293), .A2(KEYINPUT88), .B1(KEYINPUT15), .B2(new_n252), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT89), .B(G952), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  NAND2_X1  g110(.A1(G234), .A2(G237), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n292), .A2(G953), .A3(new_n297), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT21), .B(G898), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n291), .A2(new_n294), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n306));
  INV_X1    g120(.A(new_n190), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n213), .A2(new_n227), .ZN(new_n308));
  OR3_X1    g122(.A1(new_n208), .A2(KEYINPUT83), .A3(KEYINPUT19), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT83), .B1(new_n208), .B2(KEYINPUT19), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(KEYINPUT19), .B2(new_n206), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n308), .B1(new_n312), .B2(new_n215), .ZN(new_n313));
  INV_X1    g127(.A(new_n211), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n307), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n244), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G475), .A2(G902), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n306), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n317), .ZN(new_n319));
  AOI211_X1 g133(.A(KEYINPUT20), .B(new_n319), .C1(new_n244), .C2(new_n315), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n251), .B(new_n305), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n215), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n271), .A2(G146), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT0), .A4(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n202), .A2(new_n203), .ZN(new_n328));
  XNOR2_X1  g142(.A(G143), .B(G146), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT0), .B(G128), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n325), .A2(KEYINPUT1), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G128), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n325), .B(new_n326), .C1(KEYINPUT1), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n331), .B1(new_n337), .B2(new_n328), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT78), .B(G224), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n192), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n263), .A3(G104), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n189), .A2(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(G101), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(new_n342), .A3(new_n344), .A4(new_n345), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G116), .B(G119), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT2), .B(G113), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G113), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT2), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n346), .A2(new_n360), .A3(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n350), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G119), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G116), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n260), .A2(G119), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT5), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(G113), .C1(KEYINPUT5), .C2(new_n364), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n189), .A2(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n263), .A2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(G101), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n367), .A2(new_n349), .A3(new_n358), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(G110), .B(G122), .Z(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n379));
  AND4_X1   g193(.A1(new_n378), .A2(new_n372), .A3(new_n379), .A4(new_n373), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n375), .B1(new_n362), .B2(new_n371), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n381), .B2(new_n379), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n341), .B(new_n377), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT79), .B(KEYINPUT7), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n192), .B2(new_n339), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n338), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n373), .B(KEYINPUT8), .Z(new_n387));
  INV_X1    g201(.A(new_n366), .ZN(new_n388));
  OAI21_X1  g202(.A(G113), .B1(new_n364), .B2(KEYINPUT5), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n358), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n349), .A2(new_n370), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n367), .A2(new_n358), .B1(new_n349), .B2(new_n370), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n386), .A2(new_n376), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n338), .A2(KEYINPUT7), .A3(new_n340), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT80), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n338), .A2(new_n398), .A3(KEYINPUT7), .A4(new_n340), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n383), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G210), .B1(G237), .B2(G902), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n383), .A2(new_n401), .A3(new_n403), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n324), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G469), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n334), .A2(new_n336), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(KEYINPUT10), .A3(new_n349), .A4(new_n370), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n350), .A2(new_n412), .A3(new_n361), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n255), .B2(G137), .ZN(new_n415));
  INV_X1    g229(.A(G137), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT11), .A3(G134), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n255), .A2(G137), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G131), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n415), .A2(new_n417), .A3(new_n230), .A4(new_n418), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(KEYINPUT64), .A3(G131), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n349), .A2(new_n334), .A3(new_n336), .A4(new_n370), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n410), .A2(new_n413), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G110), .B(G140), .ZN(new_n430));
  INV_X1    g244(.A(G227), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G953), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n430), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n425), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n391), .A2(new_n337), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n426), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n436), .B(new_n438), .C1(KEYINPUT76), .C2(KEYINPUT12), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n423), .A2(KEYINPUT76), .A3(new_n424), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n437), .A2(new_n426), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n440), .B(new_n441), .C1(new_n442), .C2(new_n425), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n435), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n410), .A2(new_n413), .A3(new_n428), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n424), .A3(new_n423), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n434), .B1(new_n446), .B2(new_n429), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n408), .B(new_n285), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n434), .A3(new_n429), .ZN(new_n449));
  INV_X1    g263(.A(new_n429), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n439), .B2(new_n443), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(G469), .C1(new_n451), .C2(new_n434), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n408), .A2(new_n187), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n448), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G221), .ZN(new_n456));
  INV_X1    g270(.A(new_n278), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n187), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n322), .A2(new_n407), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n255), .A2(G137), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n416), .A2(G134), .ZN(new_n464));
  OAI21_X1  g278(.A(G131), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n422), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n422), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n409), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n423), .A2(new_n412), .A3(new_n424), .ZN(new_n471));
  INV_X1    g285(.A(new_n359), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n196), .A2(G210), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT27), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G101), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n474), .B(KEYINPUT27), .ZN(new_n479));
  INV_X1    g293(.A(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT67), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT30), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n423), .A2(new_n412), .A3(new_n424), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n422), .A2(new_n465), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n422), .B2(new_n465), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n489), .A2(new_n490), .A3(new_n337), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT30), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n359), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n473), .A2(new_n495), .A3(new_n483), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n485), .A2(new_n494), .A3(KEYINPUT31), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n473), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n359), .B1(new_n487), .B2(new_n491), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT28), .A4(new_n472), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n482), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT32), .ZN(new_n512));
  NOR2_X1   g326(.A1(G472), .A2(G902), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n499), .A2(new_n500), .B1(new_n506), .B2(new_n509), .ZN(new_n515));
  INV_X1    g329(.A(new_n513), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT32), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n503), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n470), .A2(new_n471), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n519), .B(new_n520), .C1(new_n472), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n522), .B2(KEYINPUT28), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n482), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT29), .B1(new_n527), .B2(new_n508), .ZN(new_n528));
  INV_X1    g342(.A(new_n494), .ZN(new_n529));
  INV_X1    g343(.A(new_n473), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n482), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n292), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n514), .A2(new_n517), .B1(G472), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n279), .B1(new_n285), .B2(G234), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n363), .B2(G128), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n363), .A2(G128), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT23), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT23), .B1(new_n335), .B2(G119), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n335), .A2(G119), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G110), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n540), .A2(new_n543), .A3(KEYINPUT73), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n539), .A2(new_n542), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT24), .B(G110), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n227), .B(new_n209), .C1(new_n547), .C2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n540), .A2(new_n543), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(G110), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n236), .B2(new_n237), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n557), .A3(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n285), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT25), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n563), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n564), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n536), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n535), .A2(G902), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT74), .B1(new_n534), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n533), .A2(G472), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n512), .B1(new_n511), .B2(new_n513), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n515), .A2(KEYINPUT32), .A3(new_n516), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n573), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n462), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n348), .ZN(G3));
  OAI21_X1  g397(.A(G472), .B1(new_n515), .B2(new_n292), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n511), .A2(new_n513), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n574), .A2(new_n460), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n211), .B1(new_n235), .B2(new_n243), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n307), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n591), .B2(new_n244), .ZN(new_n592));
  INV_X1    g406(.A(G475), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n318), .A2(new_n320), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n287), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT90), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n288), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n284), .A2(new_n595), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT91), .A4(new_n599), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n285), .A2(G478), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n605), .A2(new_n606), .B1(G478), .B2(new_n293), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n594), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n407), .A2(new_n304), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n589), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n291), .A2(new_n294), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n316), .A2(new_n317), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT20), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n316), .A2(new_n306), .A3(new_n317), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(KEYINPUT93), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT93), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n318), .B2(new_n320), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n611), .A2(new_n251), .A3(new_n617), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n589), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n558), .B(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n571), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n569), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n629), .B1(new_n586), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n407), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n321), .A2(new_n635), .A3(new_n460), .ZN(new_n636));
  INV_X1    g450(.A(new_n633), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n637), .A2(new_n584), .A3(new_n585), .A4(KEYINPUT94), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NOR3_X1   g455(.A1(new_n635), .A2(new_n460), .A3(new_n633), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(new_n579), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n299), .B1(new_n301), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n617), .B1(new_n592), .B2(new_n593), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n645), .B(new_n646), .C1(new_n621), .C2(new_n623), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT95), .B(G128), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G30));
  NAND2_X1  g464(.A1(new_n522), .A2(new_n509), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n497), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n187), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n514), .A2(new_n517), .B1(G472), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n383), .A2(new_n401), .A3(new_n403), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n403), .B1(new_n383), .B2(new_n401), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n324), .B1(new_n291), .B2(new_n294), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n594), .A2(new_n633), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n654), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n645), .B(new_n662), .Z(new_n663));
  OR2_X1    g477(.A1(new_n460), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n664), .B(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT97), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n661), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  INV_X1    g486(.A(new_n645), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n594), .A2(new_n607), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n643), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  OAI21_X1  g490(.A(new_n285), .B1(new_n444), .B2(new_n447), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(G469), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n459), .A3(new_n448), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n579), .A2(new_n573), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n612), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G15));
  NOR2_X1   g498(.A1(new_n680), .A2(new_n625), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n260), .ZN(G18));
  NAND3_X1  g500(.A1(new_n678), .A2(new_n459), .A3(new_n448), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n635), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n579), .A2(new_n322), .A3(new_n688), .A4(new_n637), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT99), .B(G119), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G21));
  OAI21_X1  g505(.A(new_n501), .B1(new_n523), .B2(new_n508), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n513), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n584), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n405), .A2(new_n406), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n594), .A2(new_n696), .A3(new_n659), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n687), .A2(new_n303), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n695), .A2(new_n697), .A3(new_n573), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G122), .ZN(G24));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n674), .A3(new_n688), .A4(new_n637), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n693), .A2(new_n637), .A3(new_n584), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n594), .A2(new_n607), .A3(new_n673), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n688), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NOR2_X1   g523(.A1(new_n534), .A2(new_n574), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT102), .B1(new_n657), .B2(new_n323), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n405), .A2(KEYINPUT102), .A3(new_n323), .A4(new_n406), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n455), .A2(KEYINPUT101), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n448), .A2(new_n452), .A3(new_n717), .A4(new_n454), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n716), .A2(new_n459), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n711), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n405), .A2(new_n323), .A3(new_n406), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n713), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n459), .A3(new_n718), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n724), .A2(KEYINPUT103), .A3(new_n725), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n710), .B(new_n674), .C1(new_n720), .C2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT42), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT103), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n719), .A2(new_n711), .A3(new_n723), .A4(new_n713), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n710), .A4(new_n674), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT104), .B(G131), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G33));
  OAI211_X1 g550(.A(new_n710), .B(new_n647), .C1(new_n720), .C2(new_n726), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  AOI22_X1  g552(.A1(new_n619), .A2(new_n620), .B1(G475), .B2(new_n250), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n607), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT43), .A3(new_n607), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(KEYINPUT105), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n587), .A2(new_n633), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n745), .A2(KEYINPUT44), .A3(new_n746), .A4(new_n747), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n449), .B1(new_n451), .B2(new_n434), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n408), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n453), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n448), .B1(new_n756), .B2(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n459), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(new_n663), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n724), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT106), .B(G137), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(KEYINPUT47), .B(new_n459), .C1(new_n757), .C2(new_n758), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n724), .A2(new_n704), .A3(new_n573), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n534), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n579), .B(new_n642), .C1(new_n647), .C2(new_n674), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n706), .B1(new_n705), .B2(new_n688), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n679), .A2(new_n407), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n703), .A2(new_n704), .A3(new_n776), .A4(KEYINPUT100), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n645), .B(KEYINPUT107), .Z(new_n780));
  NOR3_X1   g594(.A1(new_n569), .A2(new_n632), .A3(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n594), .A2(new_n781), .A3(new_n696), .A4(new_n659), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n725), .ZN(new_n783));
  INV_X1    g597(.A(new_n654), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n779), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n654), .A2(new_n782), .A3(KEYINPUT108), .A4(new_n725), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n773), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n784), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT108), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n784), .A3(new_n779), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n708), .A3(KEYINPUT52), .A4(new_n774), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n251), .B(new_n617), .C1(new_n318), .C2(new_n320), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n608), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n587), .A3(new_n611), .A4(new_n588), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n639), .A2(new_n689), .A3(new_n699), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n680), .B1(new_n625), .B2(new_n612), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n582), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n732), .A2(new_n705), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n251), .A2(new_n291), .A3(new_n294), .A4(new_n673), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n802), .A2(new_n460), .A3(new_n633), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n579), .A3(new_n715), .A4(new_n624), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n737), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n734), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n772), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(new_n793), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n737), .A2(new_n801), .A3(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n729), .B2(new_n733), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n811), .A3(KEYINPUT53), .A4(new_n800), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n807), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n734), .A2(new_n800), .A3(new_n805), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .A3(KEYINPUT53), .A4(new_n809), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n813), .B1(KEYINPUT54), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n724), .A2(new_n298), .A3(new_n687), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n744), .A2(new_n820), .A3(new_n710), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n694), .A2(new_n298), .A3(new_n574), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n744), .A2(new_n688), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n820), .A2(new_n573), .A3(new_n609), .A4(new_n654), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n822), .A2(new_n296), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n594), .A2(new_n607), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n820), .A2(new_n573), .A3(new_n654), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n744), .A2(new_n820), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n703), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n687), .A2(new_n323), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n658), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT113), .B1(new_n658), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n744), .A2(new_n823), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n658), .A2(new_n833), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n658), .A2(KEYINPUT113), .A3(new_n833), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT50), .A3(new_n744), .A4(new_n823), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n827), .B(new_n831), .C1(new_n838), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n678), .A2(new_n448), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(KEYINPUT111), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n458), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n766), .A2(new_n767), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n744), .A2(new_n854), .A3(new_n715), .A4(new_n823), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n744), .A2(new_n715), .A3(new_n823), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT110), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n766), .A2(KEYINPUT114), .A3(new_n767), .A4(new_n850), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n826), .B1(new_n845), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n857), .A3(new_n855), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT112), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n831), .B1(new_n838), .B2(new_n844), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n851), .A2(new_n857), .A3(new_n864), .A4(new_n855), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n827), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n860), .A2(new_n867), .A3(KEYINPUT115), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT115), .B1(new_n860), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n819), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(G952), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n192), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n573), .A2(new_n323), .A3(new_n459), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(KEYINPUT49), .B2(new_n846), .ZN(new_n876));
  INV_X1    g690(.A(new_n740), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n846), .A2(KEYINPUT49), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n658), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n784), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(KEYINPUT116), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n819), .A2(new_n870), .B1(new_n872), .B2(new_n192), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n880), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n192), .A2(G952), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT120), .Z(new_n888));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n377), .B1(new_n380), .B2(new_n382), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n341), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT55), .Z(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT56), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n285), .B1(new_n807), .B2(new_n812), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n889), .B(new_n896), .C1(new_n897), .C2(new_n404), .ZN(new_n898));
  INV_X1    g712(.A(new_n812), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n816), .B2(new_n809), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n404), .B(new_n292), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT119), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n888), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n892), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n403), .B(new_n285), .C1(new_n807), .C2(new_n812), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT117), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT121), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n907), .B2(KEYINPUT117), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n901), .A2(new_n905), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n892), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n888), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n889), .B1(new_n907), .B2(new_n896), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n901), .A2(KEYINPUT119), .A3(new_n895), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n910), .A2(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n807), .A2(new_n812), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n807), .A2(new_n808), .A3(new_n812), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n453), .B(KEYINPUT57), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n447), .B2(new_n444), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n897), .A2(new_n754), .A3(new_n755), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n887), .B1(new_n928), .B2(new_n929), .ZN(G54));
  AND3_X1   g744(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(new_n316), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n316), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n887), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  AOI211_X1 g750(.A(new_n605), .B(new_n936), .C1(new_n923), .C2(new_n924), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n819), .A2(new_n936), .ZN(new_n938));
  AOI211_X1 g752(.A(new_n915), .B(new_n937), .C1(new_n938), .C2(new_n605), .ZN(G63));
  XNOR2_X1  g753(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n279), .A2(new_n187), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n922), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n570), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n915), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n631), .B(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n339), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n950), .B2(new_n302), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n800), .B2(G953), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n890), .B1(G898), .B2(new_n192), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  INV_X1    g768(.A(new_n493), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n490), .A2(new_n337), .ZN(new_n956));
  INV_X1    g770(.A(new_n489), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT30), .B1(new_n958), .B2(new_n471), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(new_n312), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT124), .ZN(new_n962));
  INV_X1    g776(.A(new_n778), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n671), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n575), .A2(new_n581), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n724), .A2(new_n664), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n796), .A3(new_n967), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n762), .A2(new_n965), .A3(new_n770), .A4(new_n968), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n964), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT125), .B1(new_n964), .B2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n962), .B1(new_n973), .B2(new_n192), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n762), .A2(new_n734), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n759), .A2(new_n663), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n710), .A3(new_n697), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n737), .A2(new_n770), .A3(new_n963), .A4(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n192), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n961), .B1(G900), .B2(G953), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n431), .B2(new_n644), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n531), .A2(new_n497), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n818), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n975), .A2(new_n800), .A3(new_n978), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n985), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n529), .A2(new_n530), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n482), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n987), .B1(G952), .B2(new_n192), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n482), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n969), .A2(new_n972), .A3(new_n800), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n994), .A2(KEYINPUT126), .A3(new_n985), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT126), .B1(new_n994), .B2(new_n985), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n999), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n992), .B1(new_n998), .B2(new_n1000), .ZN(G57));
endmodule


