

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(KEYINPUT28), .ZN(n720) );
  XNOR2_X1 U554 ( .A(KEYINPUT87), .B(n780), .ZN(n519) );
  XNOR2_X1 U555 ( .A(KEYINPUT27), .B(KEYINPUT90), .ZN(n695) );
  NOR2_X1 U556 ( .A1(n747), .A2(n734), .ZN(n736) );
  XNOR2_X1 U557 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n742) );
  NOR2_X1 U558 ( .A1(G2084), .A2(n700), .ZN(n691) );
  XNOR2_X1 U559 ( .A(n743), .B(n742), .ZN(n744) );
  AND2_X1 U560 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U561 ( .A1(n803), .A2(n802), .ZN(n700) );
  AND2_X1 U562 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U563 ( .A1(n781), .A2(n519), .ZN(n782) );
  NOR2_X2 U564 ( .A1(G2104), .A2(n521), .ZN(n892) );
  AND2_X1 U565 ( .A1(n521), .A2(G2104), .ZN(n889) );
  NOR2_X1 U566 ( .A1(G651), .A2(n640), .ZN(n657) );
  NOR2_X1 U567 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U568 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U569 ( .A1(G101), .A2(n889), .ZN(n520) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n520), .Z(n524) );
  NAND2_X1 U571 ( .A1(G125), .A2(n892), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT65), .B(n522), .Z(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U575 ( .A1(n893), .A2(G113), .ZN(n527) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n525), .Z(n888) );
  NAND2_X1 U578 ( .A1(n888), .A2(G137), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U581 ( .A1(G85), .A2(n649), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  INV_X1 U583 ( .A(G651), .ZN(n532) );
  NOR2_X1 U584 ( .A1(n640), .A2(n532), .ZN(n653) );
  NAND2_X1 U585 ( .A1(G72), .A2(n653), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X2 U588 ( .A(KEYINPUT1), .B(n533), .Z(n650) );
  NAND2_X1 U589 ( .A1(G60), .A2(n650), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G47), .A2(n657), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U592 ( .A1(n537), .A2(n536), .ZN(G290) );
  XOR2_X1 U593 ( .A(G2427), .B(G2435), .Z(n539) );
  XNOR2_X1 U594 ( .A(G2454), .B(G2443), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n539), .B(n538), .ZN(n546) );
  XOR2_X1 U596 ( .A(G2451), .B(KEYINPUT101), .Z(n541) );
  XNOR2_X1 U597 ( .A(G2430), .B(G2438), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U599 ( .A(n542), .B(G2446), .Z(n544) );
  XNOR2_X1 U600 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U601 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n546), .B(n545), .ZN(n547) );
  AND2_X1 U603 ( .A1(n547), .A2(G14), .ZN(G401) );
  NAND2_X1 U604 ( .A1(G64), .A2(n650), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G52), .A2(n657), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n649), .A2(G90), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G77), .A2(n653), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(G114), .A2(n893), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G102), .A2(n889), .ZN(n556) );
  AND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U620 ( .A1(G126), .A2(n892), .ZN(n558) );
  AND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U622 ( .A1(n888), .A2(G138), .ZN(n560) );
  AND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT82), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G63), .A2(n650), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G51), .A2(n657), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U628 ( .A(KEYINPUT6), .B(n565), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n653), .A2(G76), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT74), .B(n566), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n649), .A2(G89), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT4), .B(n567), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(n570), .B(KEYINPUT5), .Z(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT75), .B(n573), .Z(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT7), .B(n574), .Z(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U641 ( .A(G223), .B(KEYINPUT68), .Z(n837) );
  NAND2_X1 U642 ( .A1(n837), .A2(G567), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U644 ( .A1(n649), .A2(G81), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G68), .A2(n653), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n580) );
  XNOR2_X1 U649 ( .A(n581), .B(n580), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G56), .A2(n650), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n582), .B(KEYINPUT69), .ZN(n583) );
  XNOR2_X1 U652 ( .A(KEYINPUT14), .B(n583), .ZN(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n657), .A2(G43), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n1006) );
  INV_X1 U656 ( .A(G860), .ZN(n609) );
  OR2_X1 U657 ( .A1(n1006), .A2(n609), .ZN(G153) );
  XNOR2_X1 U658 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G79), .A2(n653), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G54), .A2(n657), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT73), .ZN(n592) );
  NAND2_X1 U664 ( .A1(G66), .A2(n650), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n649), .A2(G92), .ZN(n593) );
  XOR2_X1 U667 ( .A(KEYINPUT72), .B(n593), .Z(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U669 ( .A(KEYINPUT15), .B(n596), .ZN(n1023) );
  INV_X1 U670 ( .A(G868), .ZN(n668) );
  NAND2_X1 U671 ( .A1(n1023), .A2(n668), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U673 ( .A1(G91), .A2(n649), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G78), .A2(n653), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G53), .A2(n657), .ZN(n601) );
  XNOR2_X1 U677 ( .A(KEYINPUT67), .B(n601), .ZN(n602) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n650), .A2(G65), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G299) );
  XNOR2_X1 U681 ( .A(KEYINPUT76), .B(n668), .ZN(n606) );
  NOR2_X1 U682 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U684 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n609), .A2(G559), .ZN(n610) );
  INV_X1 U686 ( .A(n1023), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n610), .A2(n632), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n1006), .ZN(n612) );
  XOR2_X1 U690 ( .A(KEYINPUT77), .B(n612), .Z(n615) );
  NAND2_X1 U691 ( .A1(G868), .A2(n632), .ZN(n613) );
  NOR2_X1 U692 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U694 ( .A1(n892), .A2(G123), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G111), .A2(n893), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G135), .A2(n888), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G99), .A2(n889), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n956) );
  XNOR2_X1 U702 ( .A(n956), .B(G2096), .ZN(n624) );
  INV_X1 U703 ( .A(G2100), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G93), .A2(n649), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G80), .A2(n653), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n657), .A2(G55), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT78), .B(n627), .Z(n628) );
  NOR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n650), .A2(G67), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n669) );
  NAND2_X1 U713 ( .A1(n632), .A2(G559), .ZN(n666) );
  XNOR2_X1 U714 ( .A(n1006), .B(n666), .ZN(n633) );
  NOR2_X1 U715 ( .A1(G860), .A2(n633), .ZN(n634) );
  XOR2_X1 U716 ( .A(n669), .B(n634), .Z(G145) );
  NAND2_X1 U717 ( .A1(G651), .A2(G74), .ZN(n635) );
  XOR2_X1 U718 ( .A(KEYINPUT79), .B(n635), .Z(n637) );
  NAND2_X1 U719 ( .A1(n657), .A2(G49), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT80), .B(n638), .ZN(n639) );
  NOR2_X1 U722 ( .A1(n650), .A2(n639), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n640), .A2(G87), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G88), .A2(n649), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G75), .A2(n653), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G62), .A2(n650), .ZN(n646) );
  NAND2_X1 U729 ( .A1(G50), .A2(n657), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(G166) );
  NAND2_X1 U732 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U736 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n657), .A2(G48), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(G305) );
  INV_X1 U740 ( .A(G299), .ZN(n718) );
  XNOR2_X1 U741 ( .A(n718), .B(n1006), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n660), .B(n669), .ZN(n661) );
  XNOR2_X1 U743 ( .A(KEYINPUT19), .B(n661), .ZN(n663) );
  XNOR2_X1 U744 ( .A(G288), .B(G166), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U746 ( .A(n664), .B(G290), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(G305), .ZN(n908) );
  XOR2_X1 U748 ( .A(n908), .B(n666), .Z(n667) );
  NAND2_X1 U749 ( .A1(G868), .A2(n667), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U760 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U761 ( .A1(G96), .A2(n678), .ZN(n842) );
  NAND2_X1 U762 ( .A1(n842), .A2(G2106), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U764 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U765 ( .A1(G108), .A2(n680), .ZN(n841) );
  NAND2_X1 U766 ( .A1(n841), .A2(G567), .ZN(n681) );
  NAND2_X1 U767 ( .A1(n682), .A2(n681), .ZN(n913) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT81), .B(n683), .Z(n684) );
  NOR2_X1 U770 ( .A1(n913), .A2(n684), .ZN(n840) );
  NAND2_X1 U771 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U773 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n836) );
  XOR2_X1 U774 ( .A(G1981), .B(G305), .Z(n1016) );
  NOR2_X1 U775 ( .A1(G1384), .A2(G164), .ZN(n803) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n686) );
  INV_X1 U777 ( .A(KEYINPUT84), .ZN(n685) );
  XNOR2_X1 U778 ( .A(n686), .B(n685), .ZN(n802) );
  NAND2_X1 U779 ( .A1(G8), .A2(n700), .ZN(n779) );
  NOR2_X1 U780 ( .A1(G288), .A2(G1976), .ZN(n687) );
  XNOR2_X1 U781 ( .A(n687), .B(KEYINPUT97), .ZN(n1002) );
  NOR2_X1 U782 ( .A1(n779), .A2(n1002), .ZN(n688) );
  NAND2_X1 U783 ( .A1(KEYINPUT33), .A2(n688), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n1016), .A2(n689), .ZN(n770) );
  INV_X1 U785 ( .A(KEYINPUT88), .ZN(n690) );
  NAND2_X1 U786 ( .A1(n691), .A2(n690), .ZN(n732) );
  INV_X1 U787 ( .A(n691), .ZN(n692) );
  NAND2_X1 U788 ( .A1(n692), .A2(KEYINPUT88), .ZN(n731) );
  AND2_X1 U789 ( .A1(n732), .A2(n731), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n693), .A2(G8), .ZN(n749) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n779), .ZN(n747) );
  INV_X1 U792 ( .A(n700), .ZN(n694) );
  NAND2_X1 U793 ( .A1(G2072), .A2(n694), .ZN(n696) );
  XNOR2_X1 U794 ( .A(n696), .B(n695), .ZN(n698) );
  INV_X1 U795 ( .A(G1956), .ZN(n982) );
  NOR2_X1 U796 ( .A1(n982), .A2(n694), .ZN(n697) );
  NOR2_X1 U797 ( .A1(n698), .A2(n697), .ZN(n719) );
  NAND2_X1 U798 ( .A1(n719), .A2(n718), .ZN(n717) );
  XOR2_X1 U799 ( .A(G1996), .B(KEYINPUT91), .Z(n706) );
  XNOR2_X1 U800 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n706), .A2(n707), .ZN(n699) );
  NOR2_X1 U802 ( .A1(n699), .A2(n1006), .ZN(n704) );
  NAND2_X1 U803 ( .A1(G1348), .A2(n700), .ZN(n702) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n694), .ZN(n701) );
  NAND2_X1 U805 ( .A1(n702), .A2(n701), .ZN(n713) );
  NAND2_X1 U806 ( .A1(n1023), .A2(n713), .ZN(n703) );
  NAND2_X1 U807 ( .A1(n704), .A2(n703), .ZN(n712) );
  INV_X1 U808 ( .A(G1341), .ZN(n1007) );
  NAND2_X1 U809 ( .A1(n1007), .A2(n707), .ZN(n705) );
  NAND2_X1 U810 ( .A1(n705), .A2(n700), .ZN(n710) );
  INV_X1 U811 ( .A(n706), .ZN(n925) );
  NOR2_X1 U812 ( .A1(n700), .A2(n925), .ZN(n708) );
  NAND2_X1 U813 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U814 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U815 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U816 ( .A1(n713), .A2(n1023), .ZN(n714) );
  NOR2_X1 U817 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U820 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U821 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U822 ( .A(KEYINPUT29), .B(n724), .Z(n729) );
  XOR2_X1 U823 ( .A(G2078), .B(KEYINPUT25), .Z(n725) );
  XNOR2_X1 U824 ( .A(KEYINPUT89), .B(n725), .ZN(n931) );
  NOR2_X1 U825 ( .A1(n700), .A2(n931), .ZN(n727) );
  INV_X1 U826 ( .A(G1961), .ZN(n981) );
  NOR2_X1 U827 ( .A1(n694), .A2(n981), .ZN(n726) );
  NOR2_X1 U828 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U829 ( .A1(G171), .A2(n739), .ZN(n728) );
  NAND2_X1 U830 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U831 ( .A(n730), .B(KEYINPUT92), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U833 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U834 ( .A(KEYINPUT30), .B(KEYINPUT93), .ZN(n735) );
  XNOR2_X1 U835 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U836 ( .A1(n737), .A2(G168), .ZN(n738) );
  XNOR2_X1 U837 ( .A(n738), .B(KEYINPUT94), .ZN(n741) );
  NOR2_X1 U838 ( .A1(G171), .A2(n739), .ZN(n740) );
  NOR2_X1 U839 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n750) );
  INV_X1 U841 ( .A(n750), .ZN(n746) );
  NOR2_X1 U842 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n772) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  AND2_X1 U845 ( .A1(n772), .A2(n1003), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n750), .A2(G286), .ZN(n758) );
  INV_X1 U847 ( .A(G8), .ZN(n756) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n779), .ZN(n752) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n700), .ZN(n751) );
  NOR2_X1 U850 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U851 ( .A1(n753), .A2(G303), .ZN(n754) );
  XNOR2_X1 U852 ( .A(n754), .B(KEYINPUT96), .ZN(n755) );
  OR2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U854 ( .A(n759), .B(KEYINPUT32), .ZN(n771) );
  NAND2_X1 U855 ( .A1(n760), .A2(n771), .ZN(n768) );
  INV_X1 U856 ( .A(n1003), .ZN(n764) );
  NOR2_X1 U857 ( .A1(G1971), .A2(G303), .ZN(n762) );
  INV_X1 U858 ( .A(n1002), .ZN(n761) );
  NOR2_X1 U859 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U861 ( .A1(n779), .A2(n765), .ZN(n766) );
  NOR2_X1 U862 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  NOR2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n783) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n775) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U866 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n779), .A2(n776), .ZN(n781) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U870 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U873 ( .A(KEYINPUT98), .B(n784), .ZN(n818) );
  XNOR2_X1 U874 ( .A(KEYINPUT83), .B(G1986), .ZN(n785) );
  XNOR2_X1 U875 ( .A(n785), .B(G290), .ZN(n1015) );
  NAND2_X1 U876 ( .A1(G107), .A2(n893), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G131), .A2(n888), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n892), .A2(G119), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT86), .B(n788), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n889), .A2(G95), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n882) );
  NAND2_X1 U884 ( .A1(n882), .A2(G1991), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G129), .A2(n892), .ZN(n794) );
  NAND2_X1 U886 ( .A1(G141), .A2(n888), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U888 ( .A1(n889), .A2(G105), .ZN(n795) );
  XOR2_X1 U889 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n893), .A2(G117), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n902) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n902), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n823) );
  INV_X1 U895 ( .A(n823), .ZN(n955) );
  NAND2_X1 U896 ( .A1(n1015), .A2(n955), .ZN(n806) );
  INV_X1 U897 ( .A(n802), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U899 ( .A(KEYINPUT85), .B(n805), .Z(n832) );
  NAND2_X1 U900 ( .A1(n806), .A2(n832), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G140), .A2(n888), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G104), .A2(n889), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U904 ( .A(KEYINPUT34), .B(n809), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G128), .A2(n892), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G116), .A2(n893), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U908 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U910 ( .A(KEYINPUT36), .B(n815), .Z(n905) );
  XOR2_X1 U911 ( .A(KEYINPUT37), .B(G2067), .Z(n831) );
  AND2_X1 U912 ( .A1(n905), .A2(n831), .ZN(n964) );
  NAND2_X1 U913 ( .A1(n964), .A2(n832), .ZN(n819) );
  AND2_X1 U914 ( .A1(n816), .A2(n819), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n830) );
  INV_X1 U916 ( .A(n819), .ZN(n828) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n902), .ZN(n950) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n882), .ZN(n820) );
  XOR2_X1 U920 ( .A(KEYINPUT99), .B(n820), .Z(n957) );
  NOR2_X1 U921 ( .A1(n821), .A2(n957), .ZN(n822) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n950), .A2(n824), .ZN(n825) );
  XNOR2_X1 U924 ( .A(KEYINPUT39), .B(n825), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n826), .A2(n832), .ZN(n827) );
  OR2_X1 U926 ( .A1(n828), .A2(n827), .ZN(n829) );
  AND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n834) );
  NOR2_X1 U928 ( .A1(n905), .A2(n831), .ZN(n953) );
  NAND2_X1 U929 ( .A1(n953), .A2(n832), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G188) );
  XOR2_X1 U937 ( .A(G96), .B(KEYINPUT102), .Z(G221) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n843), .B(KEYINPUT103), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U944 ( .A(G1996), .B(KEYINPUT106), .ZN(n853) );
  XOR2_X1 U945 ( .A(G1956), .B(G1961), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1991), .B(G1981), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G1966), .B(G1971), .Z(n847) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1976), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2474), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT105), .B(G2090), .Z(n857) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2678), .B(G2096), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n863) );
  XOR2_X1 U964 ( .A(G2078), .B(G2084), .Z(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n892), .ZN(n864) );
  XOR2_X1 U967 ( .A(KEYINPUT107), .B(n864), .Z(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G136), .A2(n888), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U971 ( .A(KEYINPUT108), .B(n868), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G112), .A2(n893), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G100), .A2(n889), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G130), .A2(n892), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G118), .A2(n893), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n889), .A2(G106), .ZN(n875) );
  XOR2_X1 U980 ( .A(KEYINPUT109), .B(n875), .Z(n877) );
  NAND2_X1 U981 ( .A1(n888), .A2(G142), .ZN(n876) );
  NAND2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n887) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n881) );
  XNOR2_X1 U986 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U987 ( .A(KEYINPUT110), .B(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(G164), .B(KEYINPUT111), .ZN(n884) );
  XNOR2_X1 U989 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U990 ( .A(n887), .B(n886), .Z(n900) );
  NAND2_X1 U991 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U994 ( .A1(G127), .A2(n892), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G115), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n945) );
  XNOR2_X1 U999 ( .A(G160), .B(n945), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(G162), .B(n901), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n902), .B(n956), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1006 ( .A(KEYINPUT112), .B(n908), .Z(n910) );
  XNOR2_X1 U1007 ( .A(G171), .B(G286), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(n1023), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n912), .ZN(G397) );
  INV_X1 U1011 ( .A(n913), .ZN(G319) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n916), .B(KEYINPUT114), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n919), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n920), .A2(G319), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT115), .B(n921), .Z(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1023 ( .A(G1991), .B(G25), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n930) );
  XOR2_X1 U1026 ( .A(G2067), .B(G26), .Z(n924) );
  NAND2_X1 U1027 ( .A1(n924), .A2(G28), .ZN(n928) );
  XOR2_X1 U1028 ( .A(G32), .B(n925), .Z(n926) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n926), .ZN(n927) );
  NOR2_X1 U1030 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1032 ( .A(G27), .B(n931), .Z(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT53), .B(n934), .Z(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT54), .B(G34), .Z(n935) );
  XNOR2_X1 U1036 ( .A(G2084), .B(n935), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(G35), .B(G2090), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT55), .B(n940), .ZN(n942) );
  INV_X1 U1041 ( .A(G29), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n943), .A2(G11), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(n944), .B(KEYINPUT119), .ZN(n973) );
  XOR2_X1 U1045 ( .A(G2072), .B(n945), .Z(n947) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n946) );
  NOR2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1048 ( .A(KEYINPUT50), .B(n948), .Z(n967) );
  XOR2_X1 U1049 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1051 ( .A(KEYINPUT51), .B(n951), .Z(n962) );
  XOR2_X1 U1052 ( .A(G2084), .B(G160), .Z(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1056 ( .A(KEYINPUT116), .B(n958), .Z(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT117), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT52), .B(n968), .ZN(n970) );
  INV_X1 U1063 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(G29), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1032) );
  XOR2_X1 U1067 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G1986), .B(G24), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G1971), .B(G22), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n978) );
  XOR2_X1 U1071 ( .A(G1976), .B(KEYINPUT124), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G23), .B(n976), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n980), .B(n979), .ZN(n998) );
  XNOR2_X1 U1075 ( .A(G5), .B(n981), .ZN(n996) );
  XNOR2_X1 U1076 ( .A(n982), .B(G20), .ZN(n991) );
  XOR2_X1 U1077 ( .A(G1981), .B(G6), .Z(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G4), .Z(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT123), .B(n983), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(G1348), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT122), .B(n1007), .Z(n987) );
  XNOR2_X1 U1083 ( .A(G19), .B(n987), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(n992), .B(KEYINPUT60), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G21), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1091 ( .A(KEYINPUT126), .B(n999), .Z(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT61), .ZN(n1001) );
  NOR2_X1 U1093 ( .A1(G16), .A2(n1001), .ZN(n1029) );
  XNOR2_X1 U1094 ( .A(n1002), .B(KEYINPUT120), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(n1005), .B(KEYINPUT121), .ZN(n1022) );
  XNOR2_X1 U1097 ( .A(n1007), .B(n1006), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G303), .B(G1971), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(G299), .B(G1956), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(G171), .B(G1961), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G168), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT57), .B(n1018), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XNOR2_X1 U1110 ( .A(G1348), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(G16), .B(KEYINPUT56), .Z(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(n1030), .B(KEYINPUT127), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1033), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

