//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT13), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G1gat), .B2(new_n206), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(G43gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G50gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT15), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT89), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n216), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n217), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n230), .A2(KEYINPUT15), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n227), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n229), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n213), .A2(new_n215), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(new_n217), .B2(new_n224), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n226), .B1(new_n230), .B2(KEYINPUT15), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT90), .A3(new_n239), .ZN(new_n240));
  AOI211_X1 g039(.A(KEYINPUT91), .B(new_n228), .C1(new_n235), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n240), .ZN(new_n243));
  INV_X1    g042(.A(new_n228), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n211), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n233), .A2(new_n234), .A3(new_n229), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT90), .B1(new_n238), .B2(new_n239), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT91), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n228), .B1(new_n235), .B2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n210), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n205), .B1(new_n246), .B2(new_n253), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n241), .A2(new_n245), .A3(KEYINPUT17), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n211), .B1(new_n256), .B2(new_n249), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n203), .B(new_n253), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n250), .A2(new_n256), .A3(new_n252), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n210), .B1(KEYINPUT17), .B2(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n253), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G169gat), .B(G197gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n260), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n260), .B2(new_n264), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n259), .ZN(new_n274));
  INV_X1    g073(.A(new_n254), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n264), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n270), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n264), .A3(new_n270), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(KEYINPUT92), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT22), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G211gat), .B(G218gat), .Z(new_n290));
  OR2_X1    g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n290), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n283), .B1(new_n293), .B2(KEYINPUT29), .ZN(new_n294));
  XOR2_X1   g093(.A(G141gat), .B(G148gat), .Z(new_n295));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(KEYINPUT74), .A2(new_n297), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G155gat), .B(G162gat), .Z(new_n304));
  OAI211_X1 g103(.A(new_n297), .B(new_n295), .C1(new_n304), .C2(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n294), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n283), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n293), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n308), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT31), .B(G50gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G22gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(KEYINPUT79), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n321), .B2(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT75), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT75), .B1(new_n303), .B2(new_n305), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n291), .B(KEYINPUT77), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n292), .B(KEYINPUT78), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n330), .A2(new_n313), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n314), .B(new_n323), .C1(new_n331), .C2(new_n309), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n309), .B1(new_n330), .B2(new_n313), .ZN(new_n333));
  INV_X1    g132(.A(new_n314), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n322), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT66), .ZN(new_n338));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT1), .ZN(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n343), .B(KEYINPUT66), .C1(KEYINPUT1), .C2(new_n339), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n307), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n337), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n348), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n353), .B(KEYINPUT4), .C1(new_n324), .C2(new_n325), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT3), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n310), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n307), .B2(new_n348), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n354), .A2(new_n350), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n356), .A2(new_n337), .A3(new_n350), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n353), .B(new_n357), .C1(new_n324), .C2(new_n325), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT4), .B1(new_n307), .B2(new_n348), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n364), .A3(KEYINPUT76), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(new_n361), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT0), .ZN(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT6), .ZN(new_n375));
  INV_X1    g174(.A(new_n367), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n376), .A2(new_n365), .B1(new_n359), .B2(new_n352), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(new_n372), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n368), .A2(new_n373), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(G169gat), .B2(G176gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT26), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT27), .B(G183gat), .ZN(new_n389));
  INV_X1    g188(.A(G190gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(KEYINPUT28), .A3(new_n390), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT65), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(G169gat), .B2(G176gat), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n397), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  OR3_X1    g197(.A1(new_n386), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT64), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n385), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(KEYINPUT64), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n399), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n404), .A2(new_n401), .ZN(new_n411));
  OR3_X1    g210(.A1(new_n410), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n395), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n382), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT71), .ZN(new_n415));
  INV_X1    g214(.A(new_n293), .ZN(new_n416));
  INV_X1    g215(.A(new_n395), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT25), .B1(new_n400), .B2(new_n406), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n410), .A2(new_n411), .A3(new_n408), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT70), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n417), .B(KEYINPUT70), .C1(new_n418), .C2(new_n419), .ZN(new_n423));
  INV_X1    g222(.A(new_n382), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n382), .C1(new_n413), .C2(KEYINPUT29), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n415), .A2(new_n416), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(new_n423), .A3(new_n311), .A4(new_n382), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n293), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G8gat), .B(G36gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT72), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n431), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n438), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n428), .A2(new_n431), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT30), .B1(new_n442), .B2(new_n436), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n431), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n336), .B1(new_n381), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n413), .A2(new_n348), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n420), .A2(new_n353), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(G227gat), .A4(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G15gat), .B(G43gat), .Z(new_n457));
  XNOR2_X1  g256(.A(G71gat), .B(G99gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(KEYINPUT32), .C1(new_n455), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n464));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n451), .ZN(new_n466));
  INV_X1    g265(.A(new_n452), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT69), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  AND2_X1   g271(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n465), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n460), .A2(new_n470), .A3(new_n474), .A4(new_n462), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n476), .A2(KEYINPUT36), .A3(new_n477), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n449), .A2(new_n450), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n336), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n440), .A2(new_n439), .B1(new_n443), .B2(new_n446), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(new_n380), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT80), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n428), .A2(new_n489), .A3(new_n431), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n435), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT38), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n415), .A2(new_n293), .A3(new_n425), .A4(new_n427), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n429), .A2(new_n416), .A3(new_n430), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT37), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT85), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n493), .A2(new_n497), .A3(new_n494), .A4(KEYINPUT37), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT86), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT6), .B1(new_n368), .B2(new_n373), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n377), .A2(new_n372), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n444), .A2(KEYINPUT37), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n435), .A3(new_n490), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n445), .B1(new_n510), .B2(KEYINPUT38), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(new_n506), .A3(new_n504), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n508), .A2(new_n511), .A3(new_n374), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n485), .B1(new_n503), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT82), .ZN(new_n515));
  AOI211_X1 g314(.A(KEYINPUT39), .B(new_n350), .C1(new_n364), .C2(new_n356), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT81), .B1(new_n516), .B2(new_n373), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n364), .A2(new_n356), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n351), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n518), .B(new_n372), .C1(new_n520), .C2(KEYINPUT39), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n349), .A2(new_n351), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(KEYINPUT39), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n520), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n515), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n517), .A2(new_n521), .B1(new_n520), .B2(new_n524), .ZN(new_n529));
  NOR3_X1   g328(.A1(new_n529), .A2(KEYINPUT82), .A3(KEYINPUT40), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n448), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(KEYINPUT40), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT83), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n368), .A2(new_n373), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(KEYINPUT83), .A3(KEYINPUT40), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n484), .B(new_n488), .C1(new_n514), .C2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n336), .B1(new_n476), .B2(new_n477), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(new_n380), .A3(new_n441), .A4(new_n447), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n486), .A2(new_n544), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n512), .A2(new_n374), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(new_n507), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n545), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n477), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n474), .A2(new_n470), .B1(new_n460), .B2(new_n462), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n485), .B(new_n544), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n448), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n508), .A2(new_n374), .A3(new_n512), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT87), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n543), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n282), .B1(new_n539), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G134gat), .B(G162gat), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT97), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n566), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n569), .A2(new_n573), .A3(new_n576), .A4(new_n574), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT100), .B1(new_n578), .B2(new_n579), .ZN(new_n581));
  OAI22_X1  g380(.A1(new_n249), .A2(new_n256), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n241), .A2(new_n245), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(new_n256), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n580), .A2(new_n581), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n250), .A2(new_n252), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(G190gat), .B1(new_n584), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n583), .B2(new_n585), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n578), .A2(new_n579), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n579), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT17), .A2(new_n251), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n261), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n390), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n565), .B1(new_n599), .B2(new_n287), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n589), .A2(G218gat), .A3(new_n598), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n564), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n584), .A2(new_n588), .A3(G190gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n390), .B1(new_n591), .B2(new_n597), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n287), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AND4_X1   g404(.A1(KEYINPUT98), .A2(new_n605), .A3(new_n564), .A4(new_n601), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n559), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(KEYINPUT98), .A3(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n563), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n600), .A2(new_n564), .A3(new_n601), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n558), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  OR2_X1    g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G57gat), .B(G64gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n614), .A2(new_n613), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n620), .B(KEYINPUT93), .C1(new_n616), .C2(new_n615), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n622));
  INV_X1    g421(.A(G64gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(G57gat), .ZN(new_n624));
  INV_X1    g423(.A(G57gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n624), .B(new_n626), .C1(new_n625), .C2(G64gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT20), .Z(new_n635));
  OAI21_X1  g434(.A(new_n211), .B1(new_n631), .B2(new_n630), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT96), .ZN(new_n639));
  XOR2_X1   g438(.A(G127gat), .B(G155gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G183gat), .B(G211gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n592), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n617), .A2(new_n618), .B1(new_n628), .B2(new_n627), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n650), .A2(new_n621), .A3(new_n579), .A4(new_n578), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n630), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n654), .A2(new_n594), .A3(KEYINPUT10), .A4(new_n595), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n649), .A2(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n648), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n612), .A2(new_n646), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n557), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n505), .A2(new_n506), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT102), .A3(new_n374), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT102), .B1(new_n670), .B2(new_n374), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n448), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n557), .A2(new_n668), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n681), .B2(new_n486), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n478), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n681), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n482), .A2(G15gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT105), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n690), .A2(new_n691), .B1(new_n669), .B2(new_n693), .ZN(G1326gat));
  NAND3_X1  g493(.A1(new_n557), .A2(new_n336), .A3(new_n668), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AND3_X1   g496(.A1(new_n609), .A2(new_n558), .A3(new_n610), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n558), .B1(new_n609), .B2(new_n610), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n646), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(new_n667), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n557), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n222), .A3(new_n675), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n449), .A2(new_n483), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n489), .B1(new_n428), .B2(new_n431), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT38), .B1(new_n491), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n446), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n546), .A2(new_n710), .A3(new_n507), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n492), .A2(new_n499), .A3(KEYINPUT86), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n500), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n336), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n528), .A2(new_n530), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n532), .A2(new_n533), .B1(new_n373), .B2(new_n368), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n715), .A2(new_n448), .A3(new_n536), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n707), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n548), .B1(new_n545), .B2(new_n547), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n553), .A2(KEYINPUT87), .A3(new_n554), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n542), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n612), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n539), .A2(new_n556), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n700), .A2(new_n723), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n271), .A2(new_n272), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n701), .A2(new_n728), .A3(new_n667), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n724), .A2(new_n727), .A3(new_n675), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n222), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n731), .B2(new_n730), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n706), .A2(new_n733), .ZN(G1328gat));
  NAND3_X1  g533(.A1(new_n704), .A2(new_n223), .A3(new_n448), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n724), .A2(new_n727), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n739), .A2(new_n448), .A3(new_n729), .ZN(new_n740));
  OAI221_X1 g539(.A(new_n738), .B1(new_n736), .B2(new_n735), .C1(new_n740), .C2(new_n223), .ZN(G1329gat));
  NAND3_X1  g540(.A1(new_n704), .A2(new_n214), .A3(new_n478), .ZN(new_n742));
  AND4_X1   g541(.A1(new_n482), .A2(new_n724), .A3(new_n727), .A4(new_n729), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n743), .B2(new_n214), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT47), .B1(new_n742), .B2(KEYINPUT108), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI221_X1 g545(.A(new_n742), .B1(KEYINPUT108), .B2(KEYINPUT47), .C1(new_n743), .C2(new_n214), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1330gat));
  NAND4_X1  g547(.A1(new_n557), .A2(new_n212), .A3(new_n336), .A4(new_n702), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n336), .A2(new_n724), .A3(new_n727), .A4(new_n729), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(new_n212), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT48), .B(new_n749), .C1(new_n750), .C2(new_n212), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1331gat));
  OAI211_X1 g554(.A(new_n449), .B(new_n483), .C1(new_n514), .C2(new_n538), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n556), .ZN(new_n757));
  INV_X1    g556(.A(new_n728), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n612), .A2(new_n758), .A3(new_n646), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n667), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT109), .B1(new_n759), .B2(new_n667), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n674), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n625), .ZN(G1332gat));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n486), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT49), .B(G64gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n767), .B2(new_n770), .ZN(G1333gat));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n764), .B2(new_n688), .ZN(new_n773));
  INV_X1    g572(.A(G71gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n760), .B(new_n761), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n478), .A4(new_n757), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n483), .A2(new_n774), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT110), .B1(new_n764), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n775), .A2(new_n781), .A3(new_n757), .A4(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n777), .A2(new_n783), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n764), .A2(new_n485), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g590(.A1(new_n701), .A2(new_n758), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n667), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n739), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n674), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n722), .B2(new_n793), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n757), .A2(new_n799), .A3(new_n612), .A4(new_n792), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n667), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n675), .A2(new_n571), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(G1336gat));
  NOR2_X1   g602(.A1(new_n486), .A2(G92gat), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n798), .A2(new_n667), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n724), .A2(new_n727), .A3(new_n448), .A4(new_n795), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G92gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n805), .A2(new_n807), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n810), .B1(new_n806), .B2(G92gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n805), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n796), .B2(new_n483), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n688), .A2(G99gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n801), .B2(new_n818), .ZN(G1338gat));
  NOR2_X1   g618(.A1(new_n485), .A2(G106gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n798), .A2(new_n667), .A3(new_n800), .A4(new_n820), .ZN(new_n821));
  AND4_X1   g620(.A1(new_n336), .A2(new_n724), .A3(new_n727), .A4(new_n795), .ZN(new_n822));
  INV_X1    g621(.A(G106gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT53), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n821), .B(new_n826), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1339gat));
  AOI21_X1  g627(.A(new_n203), .B1(new_n263), .B2(new_n253), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n246), .A2(new_n253), .A3(new_n205), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n269), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n269), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n832), .A2(new_n279), .A3(new_n667), .A4(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n653), .A2(new_n655), .A3(new_n648), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n653), .A2(new_n655), .A3(new_n840), .A4(new_n648), .ZN(new_n841));
  AOI211_X1 g640(.A(new_n837), .B(new_n656), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n663), .B1(new_n656), .B2(new_n837), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n836), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n841), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n666), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n835), .B1(new_n728), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n607), .A2(new_n850), .A3(new_n611), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n845), .A2(new_n666), .A3(new_n848), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n832), .A2(new_n834), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n279), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n607), .B2(new_n611), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n646), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n700), .A2(new_n701), .A3(new_n728), .A4(new_n794), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n336), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n674), .A2(new_n688), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n486), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G113gat), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n861), .A2(new_n862), .A3(new_n282), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n860), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n448), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(KEYINPUT116), .A3(new_n860), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n758), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n870), .B2(new_n862), .ZN(G1340gat));
  INV_X1    g670(.A(G120gat), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n861), .A2(new_n872), .A3(new_n794), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n869), .A2(new_n667), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n872), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n861), .B2(new_n646), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n646), .A2(G127gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n868), .B2(new_n877), .ZN(G1342gat));
  NOR2_X1   g677(.A1(new_n700), .A2(G134gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n869), .A2(new_n882), .A3(new_n879), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n861), .B2(new_n700), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n674), .A2(new_n448), .A3(new_n482), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT117), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n483), .A2(new_n486), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n674), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n336), .A2(KEYINPUT57), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n849), .B1(new_n273), .B2(new_n280), .ZN(new_n893));
  INV_X1    g692(.A(new_n835), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n611), .B(new_n607), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n271), .A2(new_n272), .A3(new_n202), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT92), .B1(new_n278), .B2(new_n279), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n853), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n835), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n700), .A2(new_n901), .A3(KEYINPUT118), .ZN(new_n902));
  INV_X1    g701(.A(new_n855), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n612), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n897), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n646), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n892), .B1(new_n906), .B2(new_n858), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n485), .B1(new_n857), .B2(new_n858), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(KEYINPUT57), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n281), .B(new_n891), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n701), .B1(new_n904), .B2(new_n851), .ZN(new_n913));
  NOR4_X1   g712(.A1(new_n612), .A2(new_n646), .A3(new_n758), .A4(new_n667), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n336), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n905), .B2(new_n646), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n892), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(KEYINPUT119), .A3(new_n281), .A4(new_n891), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n912), .A2(G141gat), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n908), .A2(new_n886), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(G141gat), .A3(new_n282), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(KEYINPUT58), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G141gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n856), .B1(new_n895), .B2(new_n896), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n701), .B1(new_n927), .B2(new_n902), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT57), .B(new_n336), .C1(new_n928), .C2(new_n914), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n929), .A2(new_n917), .B1(new_n890), .B2(new_n887), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n758), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT58), .B1(new_n931), .B2(new_n923), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n925), .A2(new_n932), .ZN(G1344gat));
  INV_X1    g732(.A(new_n922), .ZN(new_n934));
  INV_X1    g733(.A(G148gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n935), .A3(new_n667), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n915), .A2(KEYINPUT57), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n794), .B1(new_n887), .B2(new_n890), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n485), .A2(KEYINPUT57), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n701), .B1(new_n904), .B2(new_n895), .ZN(new_n941));
  NOR4_X1   g740(.A1(new_n612), .A2(new_n646), .A3(new_n281), .A4(new_n667), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT120), .A4(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(G148gat), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n946), .A2(new_n940), .B1(new_n915), .B2(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n939), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n937), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT59), .B(new_n935), .C1(new_n930), .C2(new_n667), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n936), .B1(new_n951), .B2(new_n952), .ZN(G1345gat));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n299), .A3(new_n701), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n930), .A2(new_n701), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n299), .ZN(G1346gat));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n300), .A3(new_n612), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n930), .A2(new_n612), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n300), .ZN(G1347gat));
  NAND3_X1  g758(.A1(new_n674), .A2(new_n478), .A3(new_n448), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n859), .ZN(new_n962));
  INV_X1    g761(.A(G169gat), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(new_n282), .ZN(new_n964));
  INV_X1    g763(.A(new_n960), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n859), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT121), .Z(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n758), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n964), .B1(new_n968), .B2(new_n963), .ZN(G1348gat));
  INV_X1    g768(.A(G176gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n967), .A2(new_n970), .A3(new_n667), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n962), .B2(new_n794), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  OAI21_X1  g772(.A(G183gat), .B1(new_n962), .B2(new_n646), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n701), .A2(new_n389), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n966), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n967), .A2(new_n390), .A3(new_n612), .ZN(new_n978));
  OAI21_X1  g777(.A(G190gat), .B1(new_n962), .B2(new_n700), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n982), .B(G190gat), .C1(new_n962), .C2(new_n700), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n981), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NOR3_X1   g785(.A1(new_n675), .A2(new_n486), .A3(new_n482), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n943), .B(new_n987), .C1(new_n908), .C2(new_n916), .ZN(new_n988));
  INV_X1    g787(.A(G197gat), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(new_n989), .A3(new_n282), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n908), .A2(new_n987), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(G197gat), .B1(new_n992), .B2(new_n758), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n990), .A2(new_n993), .ZN(G1352gat));
  OAI21_X1  g793(.A(G204gat), .B1(new_n988), .B2(new_n794), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n794), .A2(G204gat), .ZN(new_n996));
  AND2_X1   g795(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n997));
  NOR2_X1   g796(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n991), .A2(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n991), .A2(new_n996), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n995), .B(new_n999), .C1(new_n1000), .C2(new_n997), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1001), .B(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n992), .A2(new_n286), .A3(new_n701), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n646), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n286), .B1(new_n1005), .B2(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1007), .B1(new_n988), .B2(new_n646), .ZN(new_n1008));
  AOI21_X1  g807(.A(KEYINPUT63), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n947), .A2(KEYINPUT126), .A3(new_n701), .A4(new_n987), .ZN(new_n1010));
  AND4_X1   g809(.A1(KEYINPUT63), .A2(new_n1010), .A3(new_n1008), .A4(G211gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1004), .B1(new_n1009), .B2(new_n1011), .ZN(G1354gat));
  OAI21_X1  g811(.A(G218gat), .B1(new_n988), .B2(new_n700), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n992), .A2(new_n287), .A3(new_n612), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


