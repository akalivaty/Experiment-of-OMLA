//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  XNOR2_X1  g000(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(G137), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n188), .B(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT78), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .A4(KEYINPUT16), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT16), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT76), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(new_n201), .C1(new_n202), .C2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G128), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n211), .B(new_n213), .C1(G119), .C2(new_n212), .ZN(new_n214));
  XNOR2_X1  g028(.A(G119), .B(G128), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT24), .B(G110), .Z(new_n216));
  AOI22_X1  g030(.A1(new_n214), .A2(G110), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n214), .A2(G110), .B1(new_n215), .B2(new_n216), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(new_n199), .A3(new_n206), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n193), .A2(new_n195), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n221), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(new_n191), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n222), .B2(new_n224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  INV_X1    g044(.A(G234), .ZN(new_n231));
  OAI21_X1  g045(.A(G217), .B1(new_n231), .B2(G902), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT75), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT79), .ZN(new_n235));
  INV_X1    g049(.A(new_n225), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n227), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n225), .A2(KEYINPUT79), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n242), .A2(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  OAI22_X1  g059(.A1(new_n242), .A2(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n245), .A2(new_n246), .A3(new_n251), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n206), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G146), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n257), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n258), .A2(new_n264), .A3(KEYINPUT69), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT69), .B1(new_n258), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n253), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n259), .A3(new_n261), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n260), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n206), .A2(G143), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G128), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n206), .A2(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n268), .A2(new_n259), .A3(new_n261), .A4(KEYINPUT66), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n247), .A2(G134), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n244), .A2(G137), .ZN(new_n280));
  OAI21_X1  g094(.A(G131), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n252), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(KEYINPUT30), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n267), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n278), .A2(new_n252), .A3(new_n281), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n258), .A2(new_n264), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n250), .B2(new_n252), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g107(.A(new_n253), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n282), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n288), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n210), .A2(G116), .ZN(new_n299));
  INV_X1    g113(.A(G116), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n287), .A2(new_n298), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n267), .A2(new_n282), .A3(new_n309), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(G101), .ZN(new_n314));
  NOR2_X1   g128(.A1(G237), .A2(G953), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G210), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n314), .B(new_n316), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT31), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT31), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n311), .A2(new_n321), .A3(new_n312), .A4(new_n318), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n295), .A2(new_n310), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n312), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n256), .A2(new_n255), .A3(new_n257), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n258), .A2(new_n264), .A3(KEYINPUT69), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n330), .A2(new_n331), .B1(new_n250), .B2(new_n252), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n326), .B1(new_n332), .B2(new_n289), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n267), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n309), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n325), .B1(new_n323), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT72), .B1(new_n336), .B2(new_n318), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n323), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n317), .C1(new_n340), .C2(new_n325), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n320), .A2(new_n322), .A3(new_n337), .A4(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G472), .A2(G902), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT32), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n312), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n285), .A2(new_n286), .B1(new_n293), .B2(new_n297), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(new_n310), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT73), .B1(new_n351), .B2(new_n318), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n311), .A2(new_n312), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n317), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n336), .B2(new_n318), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n309), .B1(new_n267), .B2(new_n282), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT28), .B1(new_n349), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n339), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n227), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n227), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT74), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G472), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n241), .B1(new_n348), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G107), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(G101), .B(new_n373), .C1(new_n377), .C2(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(G107), .B1(new_n370), .B2(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n375), .B2(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n271), .A2(new_n276), .A3(new_n277), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n369), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n278), .A2(KEYINPUT82), .A3(new_n378), .A4(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n374), .A2(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n379), .A2(new_n380), .ZN(new_n397));
  OAI21_X1  g211(.A(G101), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n398), .A3(KEYINPUT4), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(G101), .C1(new_n396), .C2(new_n397), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n401), .C1(new_n265), .C2(new_n266), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n396), .A2(new_n397), .A3(G101), .ZN(new_n403));
  AOI21_X1  g217(.A(G104), .B1(new_n394), .B2(new_n395), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n404), .A2(new_n384), .A3(new_n372), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT10), .A3(new_n278), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n253), .B(KEYINPUT83), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n391), .A2(new_n402), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n406), .B2(new_n278), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT85), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n388), .A3(new_n390), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n294), .A2(KEYINPUT84), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n413), .A2(KEYINPUT12), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT12), .B1(new_n413), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G110), .B(G140), .Z(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT80), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n189), .A2(G227), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n409), .A2(new_n421), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n391), .A2(new_n402), .A3(new_n407), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n253), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G469), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT86), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n409), .B(new_n421), .C1(new_n415), .C2(new_n416), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT87), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n413), .A2(new_n414), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n413), .A2(KEYINPUT12), .A3(new_n414), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n409), .A4(new_n421), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n426), .A2(new_n409), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n422), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n432), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n429), .A3(new_n227), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n417), .A2(new_n422), .B1(new_n424), .B2(new_n426), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(G469), .C1(new_n445), .C2(G902), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n430), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  XOR2_X1   g263(.A(G110), .B(G122), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n399), .A2(new_n308), .A3(new_n307), .A4(new_n401), .ZN(new_n452));
  OAI21_X1  g266(.A(G113), .B1(new_n299), .B2(KEYINPUT5), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n378), .A2(new_n385), .A3(new_n456), .A4(new_n304), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n451), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n458), .A2(KEYINPUT6), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n452), .A2(new_n451), .A3(new_n457), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n452), .A2(KEYINPUT88), .A3(new_n451), .A4(new_n457), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n290), .A2(G125), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(G125), .B2(new_n278), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n189), .A2(G224), .ZN(new_n469));
  XOR2_X1   g283(.A(new_n468), .B(new_n469), .Z(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n278), .A2(G125), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n468), .B2(new_n475), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n453), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n455), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n406), .A2(new_n304), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n456), .A2(new_n304), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n386), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n450), .B(KEYINPUT8), .Z(new_n488));
  INV_X1    g302(.A(new_n468), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n473), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n476), .B(KEYINPUT91), .C1(new_n468), .C2(new_n475), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n479), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n462), .A2(new_n463), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n471), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G210), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n494), .A3(new_n496), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n449), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT9), .B(G234), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G221), .B1(new_n502), .B2(G902), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n447), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n370), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n189), .A3(G214), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(G143), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(G143), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n260), .A2(KEYINPUT92), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(G214), .A4(new_n315), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n251), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n514), .A3(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT94), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n205), .A2(new_n207), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT17), .A4(G131), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n516), .A2(new_n523), .A3(new_n517), .A4(new_n518), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n197), .A2(new_n199), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G146), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n220), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n511), .A2(new_n514), .A3(G131), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT18), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT18), .B2(G131), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n528), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n507), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G131), .B1(new_n511), .B2(new_n514), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n526), .B(KEYINPUT19), .ZN(new_n538));
  OAI221_X1 g352(.A(new_n205), .B1(new_n529), .B2(new_n537), .C1(G146), .C2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n535), .A2(new_n539), .A3(new_n507), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n536), .A2(G475), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n529), .A2(new_n537), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n523), .B1(new_n542), .B2(new_n517), .ZN(new_n543));
  INV_X1    g357(.A(new_n524), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n205), .A2(new_n207), .A3(new_n522), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n535), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n506), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT95), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n535), .A2(new_n539), .A3(new_n507), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n541), .A2(new_n551), .A3(new_n552), .A4(new_n227), .ZN(new_n553));
  INV_X1    g367(.A(G475), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n548), .A2(new_n554), .A3(new_n227), .A4(new_n550), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n536), .A2(KEYINPUT95), .A3(new_n540), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(KEYINPUT20), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT96), .B(G475), .Z(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n507), .A2(KEYINPUT97), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n525), .A2(new_n560), .A3(new_n535), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n525), .B2(new_n535), .ZN(new_n562));
  OR3_X1    g376(.A1(new_n561), .A2(new_n562), .A3(G902), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n553), .A2(new_n557), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(KEYINPUT100), .A2(G952), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT100), .A2(G952), .ZN(new_n567));
  AOI21_X1  g381(.A(G953), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(G234), .A2(G237), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT21), .B(G898), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(G902), .A3(G953), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n212), .B2(G143), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n212), .A2(G143), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT98), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(KEYINPUT13), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n260), .A2(G128), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n584), .C1(new_n272), .C2(new_n578), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G134), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n272), .A2(new_n580), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n244), .ZN(new_n589));
  XNOR2_X1  g403(.A(G116), .B(G122), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n377), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n375), .B2(new_n376), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT99), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n588), .B(new_n244), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n300), .A2(KEYINPUT14), .A3(G122), .ZN(new_n598));
  OAI211_X1 g412(.A(G107), .B(new_n598), .C1(new_n591), .C2(KEYINPUT14), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n593), .A3(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n586), .A2(G134), .B1(new_n593), .B2(new_n592), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n589), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n501), .A2(G217), .A3(new_n189), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n605), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n596), .A2(new_n600), .A3(new_n603), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n227), .ZN(new_n610));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(KEYINPUT15), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n610), .A2(new_n612), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n564), .A2(new_n577), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n368), .A2(new_n504), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AND2_X1   g433(.A1(new_n447), .A2(new_n503), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n342), .A2(new_n227), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n622), .A2(new_n344), .ZN(new_n623));
  INV_X1    g437(.A(new_n241), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n471), .A2(new_n496), .A3(new_n494), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n496), .B1(new_n471), .B2(new_n494), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n448), .B(new_n577), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n553), .A2(new_n557), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n563), .A2(new_n559), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n611), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n606), .A2(new_n633), .A3(new_n608), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n601), .A2(new_n602), .A3(new_n589), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n602), .B1(new_n601), .B2(new_n589), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n600), .A4(new_n607), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n605), .B(KEYINPUT101), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n604), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n635), .B1(KEYINPUT33), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n611), .A2(G902), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n632), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n631), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n628), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n625), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(new_n615), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n536), .A2(new_n540), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n552), .A3(new_n554), .A4(new_n227), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n555), .A2(KEYINPUT20), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT103), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n555), .A2(new_n661), .A3(KEYINPUT20), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n654), .B(new_n630), .C1(new_n658), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n628), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n625), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n193), .A2(new_n195), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n671), .A2(new_n223), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n223), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n239), .A3(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n234), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n504), .A2(new_n617), .A3(new_n623), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT37), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G110), .ZN(G12));
  AND3_X1   g493(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n346), .B1(new_n342), .B2(new_n343), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n365), .A2(new_n363), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n354), .B1(new_n353), .B2(new_n317), .ZN(new_n683));
  AOI211_X1 g497(.A(KEYINPUT73), .B(new_n318), .C1(new_n311), .C2(new_n312), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n682), .B1(new_n685), .B2(new_n356), .ZN(new_n686));
  INV_X1    g500(.A(G472), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n680), .A2(new_n681), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n571), .B1(new_n689), .B2(new_n575), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n664), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n504), .A2(new_n688), .A3(new_n676), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT105), .B(G128), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G30));
  XOR2_X1   g508(.A(new_n690), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n620), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n620), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n697), .A2(new_n699), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT40), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n626), .A2(new_n627), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n498), .A2(new_n499), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT38), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n449), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n317), .B1(new_n349), .B2(new_n358), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n319), .A2(G472), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(G472), .A2(G902), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n680), .B2(new_n681), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n564), .A2(new_n615), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n711), .A2(new_n675), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n701), .A2(new_n704), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n260), .ZN(G45));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n634), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n646), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n730), .A2(new_n632), .B1(new_n629), .B2(new_n630), .ZN(new_n731));
  INV_X1    g545(.A(new_n690), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n729), .A2(new_n646), .B1(new_n611), .B2(new_n610), .ZN(new_n734));
  NOR4_X1   g548(.A1(new_n734), .A2(new_n564), .A3(KEYINPUT109), .A4(new_n690), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n504), .A3(new_n688), .A4(new_n676), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G146), .ZN(G48));
  AND3_X1   g552(.A1(new_n442), .A2(new_n429), .A3(new_n227), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n429), .B1(new_n442), .B2(new_n227), .ZN(new_n740));
  INV_X1    g554(.A(new_n503), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n688), .A2(new_n650), .A3(new_n624), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT41), .B(G113), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT110), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n743), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n688), .A2(new_n665), .A3(new_n624), .A4(new_n742), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NAND2_X1  g562(.A1(new_n442), .A2(new_n227), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G469), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n500), .A2(new_n750), .A3(new_n503), .A4(new_n443), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n688), .A3(new_n617), .A4(new_n676), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  NOR2_X1   g567(.A1(new_n739), .A2(new_n740), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n503), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n500), .A2(new_n577), .A3(new_n721), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n339), .A2(new_n359), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n320), .B(new_n322), .C1(new_n757), .C2(new_n318), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n343), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n622), .A2(new_n624), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI22_X1  g576(.A1(new_n621), .A2(G472), .B1(new_n343), .B2(new_n758), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT111), .A3(new_n624), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n755), .B(new_n756), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(G122), .Z(G24));
  AND3_X1   g580(.A1(new_n622), .A2(new_n676), .A3(new_n759), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n736), .A2(new_n751), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n741), .A2(new_n449), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n498), .A2(new_n499), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n445), .B2(G902), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(new_n443), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n688), .A2(new_n624), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT109), .B1(new_n649), .B2(new_n690), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n731), .A2(new_n727), .A3(new_n732), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n770), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n368), .A2(KEYINPUT42), .A3(new_n736), .A4(new_n774), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  AND4_X1   g596(.A1(new_n688), .A2(new_n691), .A3(new_n774), .A4(new_n624), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n244), .ZN(G36));
  INV_X1    g598(.A(KEYINPUT46), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n445), .B(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n785), .B(G469), .C1(new_n787), .C2(G902), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n423), .A2(new_n427), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n445), .A2(KEYINPUT45), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(G469), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n788), .A2(new_n443), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n503), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n695), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n734), .A2(new_n631), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT43), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT43), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n734), .B2(new_n631), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n622), .A2(new_n344), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n676), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n707), .A2(new_n449), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT112), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n805), .B2(new_n806), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n798), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(new_n247), .ZN(G39));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n796), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n503), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n736), .A3(new_n808), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n348), .A2(new_n367), .A3(new_n241), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT113), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  AND2_X1   g635(.A1(new_n443), .A2(new_n773), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n690), .A2(new_n741), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n675), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT115), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n448), .B1(new_n626), .B2(new_n627), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n615), .A3(new_n564), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n443), .A2(new_n773), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n675), .A3(new_n829), .A4(new_n823), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n825), .A2(new_n720), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n737), .A2(new_n692), .A3(new_n768), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n675), .B1(new_n348), .B2(new_n367), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n504), .C1(new_n691), .C2(new_n736), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .A3(new_n768), .A4(new_n831), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n630), .B1(new_n658), .B2(new_n663), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n839), .B(new_n675), .C1(new_n348), .C2(new_n367), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n654), .A2(new_n690), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n620), .A3(new_n808), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n622), .A2(new_n676), .A3(new_n759), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n705), .A3(new_n771), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n778), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n845), .B(new_n783), .C1(new_n779), .C2(new_n780), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n564), .A2(new_n615), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n564), .B2(new_n648), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n628), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n620), .A2(new_n623), .A3(new_n849), .A4(new_n624), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n618), .A2(new_n677), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n752), .A2(new_n743), .A3(new_n747), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n765), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n838), .A2(new_n842), .A3(new_n846), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT117), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n853), .A2(new_n846), .A3(new_n842), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT53), .A4(new_n838), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n846), .A3(new_n842), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n837), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n834), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n832), .A2(new_n862), .A3(new_n833), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(KEYINPUT53), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n857), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n857), .A2(new_n855), .A3(new_n838), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n568), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n570), .B1(new_n800), .B2(new_n802), .ZN(new_n878));
  INV_X1    g692(.A(new_n764), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT111), .B1(new_n763), .B2(new_n624), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n742), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n710), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n448), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n883), .A3(KEYINPUT50), .A4(new_n878), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n754), .A2(KEYINPUT114), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n754), .A2(KEYINPUT114), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n741), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n814), .A2(new_n815), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n878), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n762), .B2(new_n764), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n809), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n720), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n624), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n754), .A2(new_n705), .A3(new_n771), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n570), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n564), .A3(new_n734), .A4(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n893), .A2(new_n899), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n767), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n888), .A2(new_n895), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT51), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n876), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n895), .A2(new_n903), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT51), .A3(new_n901), .A4(new_n888), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n368), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT48), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n898), .A2(new_n731), .A3(new_n900), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n906), .A2(new_n908), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n881), .A2(new_n826), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT118), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n868), .A2(new_n875), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n868), .A2(new_n875), .A3(new_n915), .A4(KEYINPUT119), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n889), .A2(new_n890), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT49), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n924), .A2(new_n882), .A3(new_n897), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(KEYINPUT49), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n771), .A3(new_n799), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(G75));
  AOI21_X1  g742(.A(new_n855), .B1(new_n869), .B2(new_n857), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n834), .A2(new_n837), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n861), .A2(new_n930), .A3(KEYINPUT53), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(G210), .A3(G902), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n466), .B(new_n470), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT55), .Z(new_n936));
  AND3_X1   g750(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n189), .A2(G952), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(G51));
  OAI211_X1 g754(.A(G902), .B(new_n872), .C1(new_n866), .C2(new_n855), .ZN(new_n941));
  INV_X1    g755(.A(new_n792), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT122), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n793), .A2(KEYINPUT57), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n793), .A2(KEYINPUT57), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n873), .A2(new_n874), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n932), .A2(KEYINPUT54), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n948), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n442), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n939), .B1(new_n947), .B2(new_n953), .ZN(G54));
  NAND2_X1  g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n871), .A2(G902), .A3(new_n872), .A4(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n655), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n939), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR4_X1   g773(.A1(new_n929), .A2(new_n931), .A3(new_n227), .A4(new_n955), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT123), .B1(new_n960), .B2(new_n655), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  NOR4_X1   g776(.A1(new_n941), .A2(new_n962), .A3(new_n958), .A4(new_n955), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n966), .B(new_n959), .C1(new_n961), .C2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G60));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n729), .B(new_n971), .C1(new_n950), .C2(new_n951), .ZN(new_n972));
  INV_X1    g786(.A(new_n939), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n868), .B2(new_n875), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n972), .B(new_n973), .C1(new_n729), .C2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n236), .B1(new_n873), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n978), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n932), .A2(new_n672), .A3(new_n673), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n973), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G66));
  INV_X1    g798(.A(G224), .ZN(new_n985));
  OAI21_X1  g799(.A(G953), .B1(new_n573), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n853), .B2(G953), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT125), .Z(new_n988));
  INV_X1    g802(.A(new_n466), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(G898), .B2(new_n189), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n988), .B(new_n990), .ZN(G69));
  NAND2_X1  g805(.A1(new_n701), .A2(new_n704), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n723), .A2(new_n724), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n836), .A2(new_n768), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n725), .B2(new_n995), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n819), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g815(.A(new_n848), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n368), .A2(new_n1002), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n702), .A2(new_n449), .A3(new_n707), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n1004), .B2(new_n811), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n700), .A2(new_n368), .A3(new_n808), .A4(new_n1002), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n798), .A2(new_n807), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n1006), .B(KEYINPUT126), .C1(new_n1007), .C2(new_n810), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(G953), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n350), .B(new_n538), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(KEYINPUT127), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n819), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT62), .B1(new_n994), .B2(new_n996), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n725), .A2(new_n998), .A3(new_n995), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1014), .B(new_n1009), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n189), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1018), .A2(new_n1019), .A3(new_n1011), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G900), .A2(G953), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n819), .A2(new_n811), .A3(new_n995), .ZN(new_n1022));
  INV_X1    g836(.A(new_n783), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n797), .A2(new_n368), .A3(new_n695), .A4(new_n827), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1022), .A2(new_n781), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1012), .B(new_n1021), .C1(new_n1025), .C2(G953), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1013), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1028), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1013), .A2(new_n1020), .A3(new_n1030), .A4(new_n1026), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1031), .ZN(G72));
  XOR2_X1   g846(.A(new_n714), .B(KEYINPUT63), .Z(new_n1033));
  INV_X1    g847(.A(new_n853), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1033), .B1(new_n1017), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n351), .A2(new_n317), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n939), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1033), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1038), .A2(new_n317), .A3(new_n351), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n685), .A2(new_n319), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n1033), .B(new_n1040), .C1(new_n860), .C2(new_n867), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(G57));
endmodule


