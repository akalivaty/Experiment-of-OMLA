//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n205), .B(new_n206), .ZN(G355));
  OAI21_X1  g0007(.A(G50), .B1(G58), .B2(G68), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n214), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n213), .B1(new_n224), .B2(KEYINPUT1), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g0026(.A(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n214), .B2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G13), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n229), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(G250), .B1(G257), .B2(G264), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g0034(.A1(new_n234), .A2(KEYINPUT0), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(KEYINPUT0), .ZN(new_n236));
  NOR4_X1   g0036(.A1(new_n225), .A2(new_n226), .A3(new_n235), .A4(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n216), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT66), .B(G50), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  XOR2_X1   g0053(.A(KEYINPUT8), .B(G58), .Z(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G20), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n210), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n257), .A2(new_n262), .B1(new_n255), .B2(new_n259), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n261), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  AND3_X1   g0067(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT79), .B1(G58), .B2(G68), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(new_n201), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n267), .B1(new_n270), .B2(new_n211), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT78), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n281), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n274), .A2(new_n211), .A3(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT7), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n278), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n271), .B1(new_n286), .B2(G68), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n265), .B1(new_n287), .B2(KEYINPUT16), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT16), .ZN(new_n289));
  INV_X1    g0089(.A(G68), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n285), .B2(new_n276), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n289), .B1(new_n291), .B2(new_n271), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n264), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  OAI211_X1 g0094(.A(G1), .B(G13), .C1(new_n273), .C2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(G223), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n296), .B1(G226), .B2(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G87), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n256), .B(G274), .C1(G41), .C2(G45), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n303), .B2(new_n217), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n300), .A2(new_n304), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(G169), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT18), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n286), .A2(G68), .ZN(new_n310));
  INV_X1    g0110(.A(new_n271), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT16), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(new_n261), .A3(new_n292), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n263), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT18), .ZN(new_n315));
  INV_X1    g0115(.A(new_n308), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G190), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n300), .A2(new_n304), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(G200), .B2(new_n307), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n313), .A2(new_n263), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n293), .A2(KEYINPUT17), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n274), .A2(new_n275), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G232), .A3(G1698), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(G226), .A3(new_n297), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n295), .A2(new_n302), .ZN(new_n335));
  INV_X1    g0135(.A(new_n301), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT76), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n301), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(G238), .A2(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT13), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n334), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n334), .B2(new_n340), .ZN(new_n345));
  OAI21_X1  g0145(.A(G190), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n334), .A2(new_n341), .A3(new_n340), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n334), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g0148(.A(G200), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n211), .A2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT69), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT69), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(G77), .A3(new_n354), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n290), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n261), .B1(new_n256), .B2(G20), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n258), .B2(G68), .ZN(new_n361));
  AOI22_X1  g0161(.A1(G68), .A2(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT11), .B1(new_n357), .B2(new_n261), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n346), .A2(new_n349), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(G169), .C1(new_n347), .C2(new_n348), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n334), .A2(new_n340), .ZN(new_n371));
  INV_X1    g0171(.A(new_n342), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n343), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G179), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n365), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(G232), .B(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n379));
  OAI211_X1 g0179(.A(G238), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n380));
  INV_X1    g0180(.A(G107), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n380), .C1(new_n381), .C2(new_n328), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n333), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n295), .A2(G244), .A3(new_n302), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n301), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n387), .A3(new_n301), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n359), .A2(G77), .ZN(new_n391));
  INV_X1    g0191(.A(G77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n259), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g0194(.A(KEYINPUT15), .B(G87), .Z(new_n395));
  INV_X1    g0195(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT72), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n351), .A3(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n254), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n394), .B1(new_n402), .B2(new_n261), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT73), .B1(new_n390), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n390), .A2(KEYINPUT73), .A3(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(new_n389), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G190), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n403), .ZN(new_n410));
  INV_X1    g0210(.A(G169), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n389), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(new_n412), .C1(G179), .C2(new_n389), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n327), .A2(new_n378), .A3(new_n409), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n336), .B1(new_n335), .B2(G226), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n328), .A2(new_n392), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n297), .A2(G222), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT67), .B(G223), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n297), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n328), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT68), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n333), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n415), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  OAI211_X1 g0225(.A(G190), .B(new_n415), .C1(new_n422), .C2(new_n423), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n352), .A2(new_n254), .A3(new_n354), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n265), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n258), .A2(G50), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n359), .B2(G50), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT9), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n359), .A2(G50), .ZN(new_n434));
  INV_X1    g0234(.A(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT9), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n429), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n425), .A2(new_n426), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT75), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n439), .A2(new_n426), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT75), .ZN(new_n444));
  INV_X1    g0244(.A(new_n441), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n425), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(KEYINPUT10), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n424), .A2(G179), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT70), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n429), .A2(new_n436), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n424), .B2(new_n411), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n414), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT86), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT25), .ZN(new_n458));
  AOI211_X1 g0258(.A(G107), .B(new_n258), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n256), .A2(G33), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n265), .A2(new_n258), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n381), .A3(G20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT81), .B(G116), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n273), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(new_n211), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n281), .A2(G20), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(G87), .ZN(new_n476));
  INV_X1    g0276(.A(G87), .ZN(new_n477));
  NOR4_X1   g0277(.A1(new_n281), .A2(KEYINPUT22), .A3(G20), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT24), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT24), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n473), .C1(new_n476), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n466), .B1(new_n483), .B2(new_n261), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n485));
  OAI211_X1 g0285(.A(G250), .B(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT87), .A2(G294), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT87), .A2(G294), .ZN(new_n488));
  OAI21_X1  g0288(.A(G33), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n485), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT88), .A4(new_n489), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n333), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n333), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G264), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n295), .A3(G274), .A4(new_n496), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n494), .A2(new_n505), .A3(new_n499), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(G179), .A3(new_n501), .A4(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n484), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n500), .A2(G190), .A3(new_n502), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n501), .A3(new_n506), .ZN(new_n510));
  INV_X1    g0310(.A(G200), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n508), .B1(new_n513), .B2(new_n484), .ZN(new_n514));
  OAI211_X1 g0314(.A(G244), .B(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n328), .A2(KEYINPUT4), .A3(G244), .A4(new_n297), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n328), .A2(G250), .A3(G1698), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n333), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n502), .B1(G257), .B2(new_n498), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n411), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n523), .A3(new_n305), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n266), .A2(G77), .ZN(new_n527));
  NAND2_X1  g0327(.A1(KEYINPUT6), .A2(G97), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n211), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n381), .B1(new_n285), .B2(new_n276), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n535), .A2(new_n534), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n265), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n259), .A2(new_n218), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n463), .B2(new_n218), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n525), .B(new_n526), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n524), .A2(G200), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT7), .B1(new_n281), .B2(new_n211), .ZN(new_n543));
  INV_X1    g0343(.A(new_n276), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n534), .B(G107), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n530), .A2(new_n531), .ZN(new_n546));
  INV_X1    g0346(.A(new_n529), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n549), .A3(new_n527), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n535), .A2(new_n534), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n261), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n540), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n522), .A2(new_n523), .A3(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n542), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(G116), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  OAI21_X1  g0359(.A(G33), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G244), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n561));
  OAI211_X1 g0361(.A(G238), .B(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n333), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n496), .A2(G274), .ZN(new_n565));
  OAI21_X1  g0365(.A(G250), .B1(new_n495), .B2(G1), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n333), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n511), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n319), .B(new_n567), .C1(new_n563), .C2(new_n333), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n328), .A2(new_n211), .A3(G68), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n350), .B2(new_n218), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n576), .A2(KEYINPUT82), .A3(new_n211), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT82), .B1(new_n576), .B2(new_n211), .ZN(new_n578));
  NOR3_X1   g0378(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n261), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n464), .A2(G87), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n397), .A2(new_n399), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n259), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n571), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n398), .B(new_n396), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n464), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT83), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n581), .A2(new_n588), .A3(new_n591), .A4(new_n584), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n564), .A2(G179), .A3(new_n568), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n567), .B1(new_n563), .B2(new_n333), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n411), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n541), .A2(new_n555), .A3(new_n586), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT84), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n498), .B2(G270), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT5), .A2(G41), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT5), .A2(G41), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n496), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G270), .A3(new_n295), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(KEYINPUT84), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n501), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n297), .C1(new_n279), .C2(new_n280), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT85), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT85), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n328), .A2(new_n608), .A3(G257), .A4(new_n297), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n297), .B1(new_n274), .B2(new_n275), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(G264), .B1(new_n281), .B2(G303), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n295), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(G200), .B1(new_n605), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n498), .A2(new_n598), .A3(G270), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n603), .A2(KEYINPUT84), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n502), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n618), .A3(G190), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n556), .A2(G116), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI22_X1  g0422(.A1(new_n463), .A2(new_n558), .B1(new_n258), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n471), .A2(G20), .ZN(new_n625));
  AOI21_X1  g0425(.A(G20), .B1(G33), .B2(G283), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n273), .A2(G97), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n260), .B2(new_n210), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT20), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n261), .B(new_n630), .C1(new_n622), .C2(new_n211), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n624), .B1(new_n629), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n614), .A2(new_n619), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT21), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n605), .A2(new_n613), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n633), .A2(new_n629), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n639), .B2(new_n623), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n615), .A2(new_n618), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(KEYINPUT21), .A3(G169), .A4(new_n634), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n638), .A2(G179), .A3(new_n634), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n636), .A2(new_n641), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n597), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n456), .A2(new_n514), .A3(new_n646), .ZN(G372));
  NAND2_X1  g0447(.A1(new_n376), .A2(new_n377), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n413), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n326), .A2(new_n366), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n318), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n448), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n454), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n596), .A2(new_n586), .ZN(new_n655));
  INV_X1    g0455(.A(new_n541), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n595), .A2(new_n589), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n585), .A2(new_n571), .B1(new_n595), .B2(new_n589), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n656), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n507), .A2(new_n503), .ZN(new_n665));
  INV_X1    g0465(.A(new_n484), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT90), .B1(new_n508), .B2(new_n668), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n541), .A2(new_n661), .A3(new_n555), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n666), .B2(new_n512), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n664), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n456), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n654), .B1(new_n677), .B2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n256), .A2(new_n211), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n635), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n668), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n645), .B2(new_n687), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n667), .A2(new_n686), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT91), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n514), .B1(new_n484), .B2(new_n686), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT92), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n699), .A3(new_n696), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n693), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n669), .A2(new_n685), .ZN(new_n703));
  INV_X1    g0503(.A(new_n700), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n695), .B2(new_n696), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n508), .A2(new_n686), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(G399));
  NOR2_X1   g0508(.A1(new_n232), .A2(G41), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n579), .A2(new_n558), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n709), .A2(new_n256), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n209), .B2(new_n709), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT28), .Z(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n676), .A2(new_n714), .A3(new_n686), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n655), .A2(new_n660), .A3(new_n656), .ZN(new_n716));
  INV_X1    g0516(.A(new_n661), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT26), .B1(new_n717), .B2(new_n541), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n718), .A3(new_n659), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n541), .A2(new_n661), .A3(new_n555), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n513), .B2(new_n484), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT94), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n667), .B2(new_n669), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n508), .A2(KEYINPUT94), .A3(new_n668), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n721), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT95), .B(new_n721), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n685), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n715), .B1(new_n729), .B2(new_n714), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n494), .A2(new_n505), .A3(new_n499), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n505), .B1(new_n494), .B2(new_n499), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(G200), .B1(new_n734), .B2(new_n501), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n484), .B1(new_n735), .B2(new_n509), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n646), .A2(new_n667), .A3(new_n736), .A4(new_n686), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n642), .A2(new_n305), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n522), .A2(new_n594), .A3(new_n523), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n742), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n734), .A2(new_n738), .A3(new_n744), .A4(new_n739), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n594), .A2(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n510), .A2(new_n642), .A3(new_n524), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n685), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n731), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n748), .B2(new_n685), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n691), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n730), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n713), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n229), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n256), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n709), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n690), .A2(new_n691), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n693), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n210), .B1(G20), .B2(new_n411), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n211), .A2(new_n319), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n305), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n511), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n216), .A2(new_n767), .B1(new_n769), .B2(new_n477), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n305), .A2(new_n511), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n281), .B(new_n770), .C1(G50), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n211), .B1(new_n775), .B2(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G97), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n211), .A2(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n775), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n783));
  XNOR2_X1  g0583(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n771), .A2(new_n779), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(new_n766), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n785), .A2(new_n290), .B1(new_n786), .B2(new_n392), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n768), .A2(new_n779), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n381), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n774), .A2(new_n778), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n767), .A2(new_n792), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n769), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n328), .B(new_n794), .C1(G303), .C2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n788), .ZN(new_n797));
  INV_X1    g0597(.A(new_n780), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G283), .A2(new_n797), .B1(new_n798), .B2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(new_n785), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G326), .A2(new_n773), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n487), .A2(new_n488), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n777), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n796), .A2(new_n799), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n764), .B1(new_n791), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n763), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n232), .A2(new_n328), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n495), .B2(new_n209), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n249), .B2(new_n495), .ZN(new_n814));
  NAND3_X1  g0614(.A1(G355), .A2(new_n231), .A3(new_n328), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(G116), .C2(new_n231), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n760), .B(new_n806), .C1(new_n810), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n809), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n689), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n762), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n676), .A2(new_n686), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n410), .A2(new_n685), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n406), .A2(new_n408), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n413), .B(new_n823), .C1(new_n824), .C2(new_n404), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT98), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n409), .A2(new_n827), .A3(new_n413), .A4(new_n823), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n413), .A2(new_n686), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n822), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n826), .A2(new_n828), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n675), .B1(new_n672), .B2(new_n671), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n686), .B(new_n834), .C1(new_n835), .C2(new_n663), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  INV_X1    g0638(.A(new_n753), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n760), .C1(new_n839), .C2(new_n837), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n763), .A2(new_n807), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n759), .B1(G77), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n786), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G107), .A2(new_n795), .B1(new_n847), .B2(new_n622), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n793), .B2(new_n780), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n800), .A2(KEYINPUT97), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n849), .B1(new_n853), .B2(G283), .ZN(new_n854));
  INV_X1    g0654(.A(G294), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n767), .A2(new_n855), .B1(new_n788), .B2(new_n477), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n328), .B(new_n856), .C1(G303), .C2(new_n773), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n778), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n785), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n767), .A2(new_n861), .B1(new_n786), .B2(new_n781), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n860), .B(new_n862), .C1(G137), .C2(new_n773), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n328), .B1(new_n788), .B2(new_n290), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n769), .A2(new_n202), .B1(new_n780), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(new_n867), .C1(G58), .C2(new_n777), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n863), .A2(KEYINPUT34), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n858), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n846), .B1(new_n871), .B2(new_n763), .ZN(new_n872));
  INV_X1    g0672(.A(new_n830), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n808), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n843), .A2(new_n874), .ZN(G384));
  OR2_X1    g0675(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n548), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(G116), .A3(new_n212), .A4(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT36), .Z(new_n879));
  NOR4_X1   g0679(.A1(new_n268), .A2(new_n269), .A3(new_n208), .A4(new_n392), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n880), .A2(KEYINPUT101), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n880), .A2(KEYINPUT101), .B1(new_n202), .B2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n256), .B(G13), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n730), .A2(new_n456), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n654), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n314), .A2(new_n316), .ZN(new_n887));
  INV_X1    g0687(.A(new_n683), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n314), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n889), .A3(new_n322), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n887), .A2(new_n889), .A3(new_n892), .A4(new_n322), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n314), .B(new_n888), .C1(new_n318), .C2(new_n326), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n310), .A2(new_n311), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n289), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n264), .B1(new_n900), .B2(new_n288), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT102), .B1(new_n901), .B2(new_n683), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n312), .A2(new_n261), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n287), .A2(KEYINPUT16), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n263), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT102), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n888), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n902), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n316), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n322), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n893), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n318), .B2(new_n326), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n898), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n648), .A2(new_n685), .ZN(new_n918));
  AND4_X1   g0718(.A1(new_n892), .A2(new_n887), .A3(new_n889), .A4(new_n322), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n902), .A2(new_n907), .A3(new_n322), .A4(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(KEYINPUT37), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n913), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n897), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n914), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n917), .B(new_n918), .C1(new_n916), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n377), .A2(new_n685), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n367), .A2(KEYINPUT14), .B1(new_n374), .B2(G179), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n370), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n378), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n413), .A2(new_n685), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n836), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n318), .A2(new_n683), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n925), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n886), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n737), .A2(new_n749), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT31), .ZN(new_n938));
  INV_X1    g0738(.A(new_n751), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n830), .A2(new_n929), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n915), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n750), .B2(new_n751), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n923), .B2(new_n914), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n942), .A2(KEYINPUT40), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n678), .B2(new_n752), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n898), .A2(new_n914), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT40), .B1(new_n948), .B2(new_n943), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n940), .A3(new_n941), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n456), .A3(new_n940), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n947), .A2(new_n952), .A3(G330), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n936), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n256), .B2(new_n756), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n936), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n884), .B1(new_n955), .B2(new_n956), .ZN(G367));
  NAND2_X1  g0757(.A1(new_n698), .A2(new_n700), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n656), .A2(new_n685), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n685), .B1(new_n538), .B2(new_n540), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n541), .A2(new_n555), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n703), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n541), .B1(new_n667), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n686), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n585), .A2(new_n686), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT103), .Z(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n659), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n661), .B2(new_n971), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n967), .A2(new_n968), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n701), .A2(new_n962), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT104), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n969), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n974), .A2(new_n976), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n979), .B1(new_n977), .B2(new_n980), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n709), .B(KEYINPUT41), .Z(new_n985));
  AOI21_X1  g0785(.A(new_n962), .B1(new_n706), .B2(new_n707), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n988), .B(new_n962), .C1(new_n706), .C2(new_n707), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n706), .A2(new_n707), .A3(new_n962), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n701), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n987), .A2(new_n989), .ZN(new_n996));
  INV_X1    g0796(.A(new_n992), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n991), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT106), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n702), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n958), .B(new_n703), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(new_n693), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n693), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(new_n754), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n995), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n985), .B1(new_n1006), .B2(new_n754), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n984), .B1(new_n1007), .B2(new_n758), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n810), .B1(new_n231), .B2(new_n583), .C1(new_n812), .C2(new_n244), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n853), .A2(G159), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n777), .A2(G68), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n772), .A2(new_n861), .B1(new_n767), .B2(new_n859), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n281), .B(new_n1012), .C1(G58), .C2(new_n795), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n202), .A2(new_n786), .B1(new_n788), .B2(new_n392), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G137), .B2(new_n798), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1017), .B1(new_n218), .B2(new_n788), .C1(new_n1018), .C2(new_n780), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n853), .B2(new_n803), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n281), .B1(new_n786), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G107), .B2(new_n777), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n769), .A2(new_n471), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1020), .B(new_n1023), .C1(KEYINPUT46), .C2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT107), .B(G311), .ZN(new_n1026));
  INV_X1    g0826(.A(G303), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n772), .A2(new_n1026), .B1(new_n767), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT108), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1016), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT47), .Z(new_n1031));
  OAI211_X1 g0831(.A(new_n759), .B(new_n1009), .C1(new_n1031), .C2(new_n764), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n809), .B2(new_n973), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1008), .A2(new_n1034), .ZN(G387));
  NAND2_X1  g0835(.A1(new_n1004), .A2(new_n709), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n754), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1036), .A2(KEYINPUT111), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(KEYINPUT111), .B2(new_n1036), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(new_n757), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n328), .B1(new_n798), .B2(G326), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n471), .B2(new_n788), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n767), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G322), .A2(new_n773), .B1(new_n1044), .B2(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n1027), .B2(new_n786), .C1(new_n852), .C2(new_n1026), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n795), .A2(new_n803), .B1(new_n777), .B2(G283), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n772), .A2(new_n781), .B1(new_n769), .B2(new_n392), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n281), .B(new_n1055), .C1(G97), .C2(new_n797), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n587), .A2(new_n777), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G50), .A2(new_n1044), .B1(new_n798), .B2(G150), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n254), .A2(new_n800), .B1(new_n847), .B2(G68), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n764), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n241), .A2(new_n495), .A3(new_n328), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n255), .B2(G50), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n710), .B1(new_n1066), .B2(new_n281), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n231), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n809), .B(new_n763), .C1(new_n232), .C2(G107), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n760), .B(new_n1061), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n958), .B2(new_n818), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT110), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1041), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1040), .A2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n709), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n990), .A2(new_n702), .A3(new_n993), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n701), .B1(new_n996), .B2(new_n998), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1078), .B2(new_n1004), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n1006), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1076), .A2(new_n1077), .A3(new_n758), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n810), .B1(new_n218), .B2(new_n231), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n252), .B2(new_n811), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n760), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT112), .Z(new_n1085));
  NAND2_X1  g0885(.A1(new_n853), .A2(G50), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n328), .B1(new_n788), .B2(new_n477), .C1(new_n255), .C2(new_n786), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G77), .B2(new_n777), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n769), .A2(new_n290), .B1(new_n780), .B2(new_n861), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT113), .Z(new_n1090));
  OAI22_X1  g0890(.A1(new_n772), .A2(new_n859), .B1(new_n767), .B2(new_n781), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n853), .A2(G303), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n772), .A2(new_n1018), .B1(new_n767), .B2(new_n793), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n769), .A2(new_n1021), .B1(new_n780), .B2(new_n792), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G294), .B2(new_n847), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n328), .B(new_n789), .C1(new_n622), .C2(new_n777), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1093), .A2(new_n1100), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1085), .B1(new_n764), .B2(new_n1101), .C1(new_n962), .C2(new_n818), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1081), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1080), .A2(new_n1103), .ZN(G390));
  AND3_X1   g0904(.A1(new_n923), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT39), .B1(new_n898), .B2(new_n914), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n932), .A2(new_n918), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n719), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT94), .B1(new_n508), .B2(new_n668), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n667), .A2(new_n669), .A3(new_n722), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n675), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1111), .B2(KEYINPUT95), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n728), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n686), .B(new_n834), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n929), .B1(new_n1114), .B2(new_n931), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n915), .B1(new_n648), .B2(new_n685), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n940), .A2(KEYINPUT114), .A3(G330), .A4(new_n941), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n941), .B(G330), .C1(new_n750), .C2(new_n751), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1107), .B(new_n1119), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n758), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT115), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT115), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1124), .A2(new_n1128), .A3(new_n758), .A4(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1116), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n930), .B1(new_n729), .B2(new_n834), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n929), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1122), .B1(new_n1133), .B2(new_n1107), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1125), .ZN(new_n1135));
  OAI211_X1 g0935(.A(G330), .B(new_n873), .C1(new_n750), .C2(new_n751), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n929), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n836), .A2(new_n931), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n753), .A2(new_n941), .B1(new_n929), .B2(new_n1136), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1140), .A2(new_n1141), .B1(new_n1132), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n456), .B(G330), .C1(new_n750), .C2(new_n751), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n885), .A2(new_n654), .A3(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n1134), .A2(new_n1135), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1144), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n653), .B(new_n1147), .C1(new_n730), .C2(new_n456), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1137), .A2(new_n1114), .A3(new_n931), .A4(new_n1119), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1118), .A2(new_n1121), .B1(new_n929), .B2(new_n1136), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1141), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1124), .A2(new_n1148), .A3(new_n1152), .A4(new_n1125), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1146), .A2(new_n709), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n808), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n281), .B1(new_n798), .B2(G125), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n781), .B2(new_n776), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n772), .A2(new_n1159), .B1(new_n767), .B2(new_n866), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n202), .A2(new_n788), .B1(new_n786), .B2(new_n1161), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1158), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT53), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n769), .B2(new_n859), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n795), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n853), .A2(G137), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G283), .A2(new_n773), .B1(new_n847), .B2(G97), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n558), .B2(new_n767), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n853), .B2(G107), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n281), .B1(new_n769), .B2(new_n477), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n788), .A2(new_n290), .B1(new_n780), .B2(new_n855), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(G77), .C2(new_n777), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1163), .A2(new_n1167), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n759), .B1(new_n254), .B2(new_n845), .C1(new_n1174), .C2(new_n764), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1156), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AND4_X1   g0977(.A1(KEYINPUT116), .A2(new_n1130), .A3(new_n1154), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1152), .A2(new_n1148), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1075), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1176), .B1(new_n1181), .B2(new_n1153), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT116), .B1(new_n1182), .B2(new_n1130), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1178), .A2(new_n1183), .ZN(G378));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n452), .A2(new_n683), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n448), .A2(new_n454), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n448), .B2(new_n454), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1186), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n455), .A2(new_n1187), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n448), .A2(new_n454), .A3(new_n1188), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n1193), .A3(new_n1185), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n951), .B2(G330), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n691), .B(new_n1195), .C1(new_n949), .C2(new_n950), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n935), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1195), .B1(new_n946), .B2(new_n691), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n925), .A2(new_n933), .A3(new_n934), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n951), .A2(G330), .A3(new_n1196), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT119), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1199), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1201), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT119), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1207), .A3(new_n758), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n760), .B1(new_n202), .B2(new_n844), .ZN(new_n1209));
  AOI211_X1 g1009(.A(G41), .B(new_n328), .C1(new_n795), .C2(G77), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n216), .B2(new_n788), .C1(new_n1021), .C2(new_n780), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT117), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G116), .A2(new_n773), .B1(new_n800), .B2(G97), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n1011), .C1(new_n381), .C2(new_n767), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n587), .B2(new_n847), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT118), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G50), .B1(new_n275), .B2(new_n294), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G125), .A2(new_n773), .B1(new_n800), .B2(G132), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n859), .B2(new_n776), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n847), .A2(G137), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n1159), .B2(new_n767), .C1(new_n769), .C2(new_n1161), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1221), .A2(new_n1223), .A3(KEYINPUT59), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n781), .B2(new_n788), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT59), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1219), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1218), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(KEYINPUT58), .B2(new_n1217), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1209), .B1(new_n1231), .B2(new_n764), .C1(new_n1196), .C2(new_n808), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1208), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1153), .A2(new_n1148), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1207), .A3(new_n1205), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1075), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G375));
  AOI22_X1  g1041(.A1(G132), .A2(new_n773), .B1(new_n1044), .B2(G137), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n852), .B2(new_n1161), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(KEYINPUT121), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n769), .A2(new_n781), .B1(new_n786), .B2(new_n859), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n328), .B1(new_n776), .B2(new_n202), .C1(new_n216), .C2(new_n788), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(G128), .C2(new_n798), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(KEYINPUT121), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n853), .A2(new_n622), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n218), .A2(new_n769), .B1(new_n767), .B2(new_n1021), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G303), .B2(new_n798), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n772), .A2(new_n855), .B1(new_n786), .B2(new_n381), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n328), .B(new_n1253), .C1(G77), .C2(new_n797), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1057), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1249), .A2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n759), .B1(G68), .B2(new_n845), .C1(new_n1256), .C2(new_n764), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n929), .B2(new_n807), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1152), .B2(new_n758), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n985), .B(KEYINPUT120), .Z(new_n1260));
  NAND2_X1  g1060(.A1(new_n1180), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1152), .A2(new_n1148), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(G381));
  NOR2_X1   g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1265), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1266));
  INV_X1    g1066(.A(G387), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1130), .A2(new_n1154), .A3(new_n1177), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .A4(new_n1240), .ZN(G407));
  INV_X1    g1070(.A(G213), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(G343), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1240), .A2(new_n1269), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(G213), .A3(new_n1273), .ZN(G409));
  AND2_X1   g1074(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1232), .B1(new_n1275), .B2(new_n757), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1234), .A2(new_n1205), .A3(new_n1207), .A4(new_n1260), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1276), .B1(new_n1278), .B2(KEYINPUT123), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1268), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT116), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1268), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1182), .A2(KEYINPUT116), .A3(new_n1130), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1240), .A2(KEYINPUT122), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT122), .B1(G378), .B2(new_n1240), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1272), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1233), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1285), .A3(new_n1286), .A4(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT122), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1282), .B1(new_n1298), .B2(new_n1287), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1299), .B2(new_n1272), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1272), .A2(G2897), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1180), .A2(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1262), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n709), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n1262), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1259), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n843), .A3(new_n874), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1259), .C1(new_n1306), .C2(new_n1305), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT124), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1302), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1310), .B(new_n1311), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1302), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT61), .B1(new_n1301), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1293), .A2(new_n1300), .A3(new_n1317), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1290), .A2(new_n1292), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1316), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1315), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n820), .B1(new_n1040), .B2(new_n1073), .ZN(new_n1324));
  OR2_X1    g1124(.A1(new_n1264), .A2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1005), .B1(new_n999), .B2(new_n702), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n701), .B1(new_n994), .B2(KEYINPUT106), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n754), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n985), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n758), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n984), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1034), .B(G390), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(G390), .B1(new_n1008), .B2(new_n1034), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1325), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(G390), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(G387), .A2(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1264), .A2(new_n1324), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1338), .A3(new_n1332), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1335), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1323), .A2(new_n1340), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1293), .A2(new_n1300), .A3(KEYINPUT63), .A4(new_n1319), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1340), .A2(KEYINPUT61), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1344), .B1(new_n1314), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1320), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1342), .B(new_n1343), .C1(new_n1346), .C2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1341), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(new_n1298), .A2(new_n1287), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1269), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  AOI22_X1  g1152(.A1(new_n1350), .A2(new_n1351), .B1(new_n1352), .B2(new_n1310), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1310), .B(KEYINPUT126), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1340), .B(new_n1354), .C1(new_n1355), .C2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1356), .A2(new_n1355), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1360), .A2(new_n1353), .ZN(new_n1361));
  OR2_X1    g1161(.A1(new_n1361), .A2(new_n1340), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1361), .A2(KEYINPUT127), .A3(new_n1340), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1359), .A2(new_n1362), .A3(new_n1363), .ZN(G402));
endmodule


