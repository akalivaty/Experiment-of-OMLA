//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n543,
    new_n544, new_n545, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1141, new_n1142,
    new_n1143, new_n1144;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n462), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT65), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT66), .Z(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(G2105), .ZN(new_n484));
  MUX2_X1   g059(.A(G100), .B(G112), .S(G2105), .Z(new_n485));
  AOI22_X1  g060(.A1(new_n484), .A2(G124), .B1(G2104), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n483), .A2(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n478), .B2(new_n462), .ZN(new_n489));
  AND2_X1   g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n472), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n478), .B2(new_n462), .ZN(new_n493));
  AND2_X1   g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n472), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT67), .A2(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(new_n501), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(new_n502), .B2(new_n503), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G166));
  XOR2_X1   g092(.A(KEYINPUT68), .B(KEYINPUT7), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n509), .A2(G89), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(new_n504), .A2(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n510), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n515), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n528), .A2(new_n530), .ZN(G171));
  NAND2_X1  g106(.A1(G68), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(G56), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n515), .B1(new_n535), .B2(KEYINPUT69), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(KEYINPUT69), .B2(new_n535), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G81), .B1(new_n504), .B2(G43), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT70), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n539), .A3(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT71), .ZN(G188));
  NAND2_X1  g121(.A1(new_n504), .A2(G53), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n515), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n509), .A2(G91), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(G299));
  INV_X1    g127(.A(G171), .ZN(G301));
  INV_X1    g128(.A(G168), .ZN(G286));
  INV_X1    g129(.A(G166), .ZN(G303));
  NAND2_X1  g130(.A1(new_n509), .A2(G87), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n504), .A2(G49), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(G288));
  INV_X1    g134(.A(G61), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n507), .B2(new_n508), .ZN(new_n561));
  AND2_X1   g136(.A1(G73), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT72), .B(G651), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n509), .A2(G86), .B1(new_n504), .B2(G48), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G305));
  NAND2_X1  g143(.A1(new_n504), .A2(G47), .ZN(new_n569));
  INV_X1    g144(.A(G85), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n510), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n515), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G301), .A2(G868), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n509), .A2(G92), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G66), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n533), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G54), .B2(new_n504), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT74), .Z(new_n585));
  OAI21_X1  g160(.A(new_n576), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n576), .B1(new_n585), .B2(G868), .ZN(G321));
  NOR2_X1   g162(.A1(G299), .A2(G868), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g164(.A(new_n588), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n591), .B2(G860), .ZN(G148));
  NAND2_X1  g167(.A1(new_n537), .A2(new_n539), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n585), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n585), .A2(new_n596), .A3(new_n591), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  MUX2_X1   g173(.A(new_n593), .B(new_n598), .S(G868), .Z(G323));
  XNOR2_X1  g174(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g175(.A(G111), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n601), .A2(KEYINPUT77), .A3(G2105), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT77), .B1(new_n601), .B2(G2105), .ZN(new_n603));
  OAI21_X1  g178(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n481), .A2(G135), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT76), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n484), .A2(new_n607), .A3(G123), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n484), .B2(G123), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(G2096), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(G2096), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2100), .Z(new_n616));
  NAND3_X1  g191(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(G156));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT15), .B(G2435), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2427), .ZN(new_n621));
  INV_X1    g196(.A(G2430), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n621), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XNOR2_X1  g209(.A(G2072), .B(G2078), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT17), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(KEYINPUT78), .ZN(new_n640));
  AOI211_X1 g215(.A(new_n634), .B(new_n639), .C1(new_n638), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT79), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n638), .A3(new_n634), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n634), .A2(new_n637), .A3(new_n635), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT18), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1956), .B(G2474), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1961), .B(G1966), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n653), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT20), .Z(new_n657));
  AOI211_X1 g232(.A(new_n655), .B(new_n657), .C1(new_n650), .C2(new_n654), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1981), .B(G1986), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G229));
  INV_X1    g240(.A(G29), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(G32), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n481), .A2(G141), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  NAND3_X1  g244(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT26), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n672));
  AOI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n484), .C2(G129), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n667), .B1(new_n674), .B2(G29), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT27), .B(G1996), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT90), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NOR2_X1   g254(.A1(G168), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n679), .B2(G21), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT91), .B(G1966), .ZN(new_n682));
  OAI22_X1  g257(.A1(new_n681), .A2(new_n682), .B1(new_n610), .B2(new_n666), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(G5), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G171), .B2(new_n679), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G1961), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G11), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT30), .B(G28), .Z(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n688), .C1(G29), .C2(new_n689), .ZN(new_n690));
  OR3_X1    g265(.A1(new_n683), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n678), .B1(KEYINPUT92), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(KEYINPUT92), .ZN(new_n693));
  NOR2_X1   g268(.A1(G29), .A2(G33), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT25), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n472), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n481), .B2(G139), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(G29), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G2072), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n675), .A2(new_n676), .ZN(new_n703));
  AND2_X1   g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  NOR2_X1   g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n666), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT88), .Z(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n474), .B2(new_n666), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G2084), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G1961), .B2(new_n686), .ZN(new_n710));
  NOR2_X1   g285(.A1(G27), .A2(G29), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G164), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2078), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n703), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n693), .A2(new_n702), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n692), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT93), .Z(new_n717));
  NOR2_X1   g292(.A1(G16), .A2(G23), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT82), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G288), .B2(new_n679), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT83), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT33), .B(G1976), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G6), .B(G305), .S(G16), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G22), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G166), .B2(G16), .ZN(new_n728));
  INV_X1    g303(.A(G1971), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n723), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT84), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT34), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n679), .A2(G24), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n574), .B(KEYINPUT81), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n679), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1986), .ZN(new_n739));
  NOR2_X1   g314(.A1(G25), .A2(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n484), .A2(G119), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n481), .A2(G131), .ZN(new_n742));
  MUX2_X1   g317(.A(G95), .B(G107), .S(G2105), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2104), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT80), .Z(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  XOR2_X1   g324(.A(new_n748), .B(new_n749), .Z(new_n750));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n739), .B(new_n750), .C1(new_n751), .C2(KEYINPUT36), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n734), .A2(new_n735), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G35), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G162), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2090), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n679), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n766));
  MUX2_X1   g341(.A(G19), .B(new_n593), .S(G16), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1341), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n666), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  MUX2_X1   g345(.A(G104), .B(G116), .S(G2105), .Z(new_n771));
  AOI22_X1  g346(.A1(new_n484), .A2(G128), .B1(G2104), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n481), .A2(G140), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n679), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n585), .B2(new_n679), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT86), .B(G1348), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n778), .B(new_n782), .C1(new_n758), .C2(G2090), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n765), .A2(new_n766), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n717), .A2(new_n755), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n753), .A2(new_n754), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n785), .A2(new_n787), .ZN(G311));
  OR2_X1    g363(.A1(new_n785), .A2(new_n787), .ZN(G150));
  XOR2_X1   g364(.A(KEYINPUT96), .B(G860), .Z(new_n790));
  AOI22_X1  g365(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n515), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n509), .A2(G93), .B1(new_n504), .B2(G55), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT37), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n794), .A2(new_n795), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n593), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n593), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT38), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n585), .A2(G559), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT39), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n790), .B1(new_n806), .B2(KEYINPUT39), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n797), .B1(new_n807), .B2(new_n808), .ZN(G145));
  XNOR2_X1  g384(.A(new_n610), .B(G160), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G162), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n746), .B(new_n614), .ZN(new_n813));
  MUX2_X1   g388(.A(G106), .B(G118), .S(G2105), .Z(new_n814));
  AOI22_X1  g389(.A1(new_n484), .A2(G130), .B1(G2104), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n481), .A2(KEYINPUT99), .A3(G142), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT99), .B1(new_n481), .B2(G142), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n813), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n674), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n700), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n774), .B(G164), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n825), .A2(new_n819), .A3(new_n826), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n812), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n827), .A2(new_n812), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n834), .B2(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g412(.A(G166), .B(G305), .Z(new_n838));
  INV_X1    g413(.A(G288), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n574), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT42), .Z(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  INV_X1    g418(.A(G299), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n584), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n584), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G299), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n584), .A3(KEYINPUT102), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(KEYINPUT41), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n845), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(KEYINPUT41), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n595), .A2(new_n597), .A3(new_n802), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n802), .B1(new_n595), .B2(new_n597), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n843), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n853), .B(KEYINPUT101), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n843), .B1(new_n858), .B2(new_n854), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n842), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n860), .A2(new_n861), .A3(new_n842), .ZN(new_n865));
  OAI211_X1 g440(.A(KEYINPUT104), .B(new_n842), .C1(new_n860), .C2(new_n861), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  MUX2_X1   g442(.A(new_n798), .B(new_n867), .S(G868), .Z(G295));
  MUX2_X1   g443(.A(new_n798), .B(new_n867), .S(G868), .Z(G331));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n871));
  NAND2_X1  g446(.A1(G301), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(G171), .A2(KEYINPUT105), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(G168), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(G286), .A2(new_n871), .A3(G301), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n801), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n799), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n802), .A2(new_n880), .A3(new_n876), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n800), .A2(new_n801), .A3(new_n874), .A4(new_n875), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n854), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n878), .A3(new_n853), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n841), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n885), .ZN(new_n889));
  INV_X1    g464(.A(new_n841), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(KEYINPUT43), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n886), .A2(new_n887), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n883), .A2(new_n859), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n882), .A2(new_n878), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n851), .A2(KEYINPUT41), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n897), .C1(KEYINPUT41), .C2(new_n853), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n841), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n893), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT44), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n888), .A2(new_n893), .A3(new_n891), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n894), .B2(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT44), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n870), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n909), .A2(new_n901), .A3(KEYINPUT107), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(G397));
  INV_X1    g486(.A(G1384), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n499), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n468), .A2(new_n473), .A3(G40), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G1996), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n820), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n774), .A2(G2067), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n772), .A2(new_n776), .A3(new_n773), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n674), .A2(G1996), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n746), .B(new_n749), .Z(new_n925));
  OAI21_X1  g500(.A(new_n917), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1986), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n574), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n917), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n930), .B(KEYINPUT108), .Z(new_n931));
  INV_X1    g506(.A(KEYINPUT54), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n913), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n499), .A2(KEYINPUT109), .A3(new_n912), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n916), .B1(new_n913), .B2(KEYINPUT50), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1961), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n941));
  INV_X1    g516(.A(G2078), .ZN(new_n942));
  INV_X1    g517(.A(new_n916), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n912), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n915), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n939), .A2(new_n940), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n499), .A2(KEYINPUT109), .A3(new_n912), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT109), .B1(new_n499), .B2(new_n912), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n914), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n499), .A2(new_n950), .A3(KEYINPUT45), .A4(new_n912), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n916), .B1(new_n944), .B2(KEYINPUT114), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n941), .A2(G2078), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n949), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G301), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT50), .ZN(new_n956));
  INV_X1    g531(.A(new_n938), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n940), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n945), .A2(new_n941), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT53), .A3(new_n942), .A4(new_n944), .ZN(new_n961));
  AND4_X1   g536(.A1(G301), .A2(new_n958), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n932), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n958), .A2(new_n954), .A3(new_n959), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G171), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n946), .A2(G301), .A3(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(KEYINPUT124), .A3(new_n932), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(G166), .B2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT55), .B(G8), .C1(new_n512), .C2(new_n516), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n943), .B1(new_n913), .B2(KEYINPUT50), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2090), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n960), .A2(new_n944), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n980), .B1(new_n729), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n934), .A2(new_n943), .A3(new_n936), .ZN(new_n985));
  INV_X1    g560(.A(new_n983), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n839), .A2(G1976), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n567), .A2(new_n563), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G1981), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(G305), .B2(G1981), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT49), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(KEYINPUT112), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n995));
  OAI221_X1 g570(.A(new_n991), .B1(new_n995), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n994), .A2(new_n986), .A3(new_n985), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n985), .A2(new_n999), .A3(new_n986), .A4(new_n987), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n989), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n975), .B(KEYINPUT110), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n937), .A2(new_n980), .A3(new_n938), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n981), .A2(new_n729), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n972), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n984), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G171), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n946), .A2(G301), .A3(new_n954), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT54), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n965), .A2(new_n970), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G168), .A2(new_n983), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(KEYINPUT51), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n952), .A2(new_n951), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n934), .B2(new_n936), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n682), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n937), .A2(new_n1020), .A3(new_n938), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n983), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1016), .B1(new_n1022), .B2(KEYINPUT123), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(KEYINPUT123), .B2(new_n1022), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n972), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT51), .B1(new_n1025), .B2(new_n1014), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1024), .A2(new_n1026), .B1(new_n1014), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT125), .B1(new_n1013), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1012), .A2(new_n1002), .A3(new_n1007), .A4(new_n984), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT124), .B1(new_n969), .B2(new_n932), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(KEYINPUT123), .A3(new_n986), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1015), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1022), .A2(KEYINPUT123), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1027), .A2(new_n1014), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT125), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1032), .A2(new_n1038), .A3(new_n1039), .A4(new_n970), .ZN(new_n1040));
  XNOR2_X1  g615(.A(G299), .B(KEYINPUT57), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT50), .B1(new_n947), .B2(new_n948), .ZN(new_n1042));
  INV_X1    g617(.A(new_n913), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n916), .B1(new_n1043), .B2(new_n935), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1956), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT118), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n960), .A2(new_n944), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1045), .A2(new_n1049), .A3(KEYINPUT119), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n1051));
  INV_X1    g626(.A(G1956), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n977), .B2(new_n978), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1053), .B2(new_n1048), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1041), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n781), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n937), .B2(new_n938), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n985), .A2(G2067), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n848), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1041), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1053), .A3(new_n1048), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NOR4_X1   g638(.A1(new_n1057), .A2(new_n1058), .A3(KEYINPUT60), .A4(new_n584), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n1057), .A2(new_n1058), .A3(new_n848), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1059), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(KEYINPUT60), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1055), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1041), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT61), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1062), .C2(new_n1069), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1067), .B(new_n1068), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n915), .A2(new_n918), .A3(new_n943), .A4(new_n944), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n960), .A2(KEYINPUT120), .A3(new_n918), .A4(new_n944), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  AOI22_X1  g655(.A1(new_n1078), .A2(new_n1079), .B1(new_n985), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1081), .B2(new_n593), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1075), .A3(new_n593), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1075), .B(KEYINPUT59), .C1(new_n1081), .C2(new_n593), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1063), .B1(new_n1074), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1029), .A2(new_n1040), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1006), .A2(new_n975), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1001), .A2(KEYINPUT113), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT113), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n989), .A2(new_n997), .A3(new_n1092), .A4(new_n1000), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT117), .B(new_n1090), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT63), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1022), .A2(KEYINPUT115), .A3(G168), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT115), .B1(new_n1022), .B2(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n1101), .B2(new_n1090), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n984), .A2(new_n1002), .A3(new_n1007), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1095), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT116), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1108), .B(new_n1095), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1101), .A2(new_n1007), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n997), .A2(new_n998), .A3(new_n839), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(G1981), .B2(G305), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(new_n986), .A3(new_n985), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1089), .A2(KEYINPUT126), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n955), .A3(new_n1008), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1100), .A2(new_n1102), .B1(new_n1106), .B2(KEYINPUT116), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1115), .B1(new_n1122), .B2(new_n1109), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT126), .B1(new_n1123), .B2(new_n1089), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n931), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n747), .A2(new_n749), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n921), .B1(new_n924), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n917), .A2(new_n927), .A3(new_n574), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT48), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n917), .A2(new_n1127), .B1(new_n926), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n922), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n917), .B1(new_n1131), .B2(new_n674), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n917), .A2(new_n918), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT46), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT47), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT127), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1125), .A2(new_n1138), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g714(.A(new_n892), .ZN(new_n1141));
  INV_X1    g715(.A(new_n900), .ZN(new_n1142));
  NOR2_X1   g716(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR4_X1   g717(.A1(G227), .A2(G229), .A3(new_n459), .A4(G401), .ZN(new_n1144));
  NAND3_X1  g718(.A1(new_n836), .A2(new_n1143), .A3(new_n1144), .ZN(G225));
  INV_X1    g719(.A(G225), .ZN(G308));
endmodule


