//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT92), .B(G8gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206));
  INV_X1    g005(.A(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(KEYINPUT91), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n204), .A2(KEYINPUT90), .A3(new_n208), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n213), .A2(G8gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n209), .B(new_n215), .C1(G1gat), .C2(new_n204), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(KEYINPUT89), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n223));
  INV_X1    g022(.A(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(G36gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT14), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n220), .A2(new_n222), .A3(new_n223), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232));
  INV_X1    g031(.A(new_n221), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT87), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT87), .ZN(new_n236));
  AOI211_X1 g035(.A(new_n232), .B(new_n223), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n234), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n236), .A3(new_n221), .ZN(new_n239));
  INV_X1    g038(.A(new_n223), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT88), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n231), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n218), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n231), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT87), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT87), .B1(new_n226), .B2(new_n228), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n246), .A2(new_n247), .A3(new_n233), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n232), .B1(new_n248), .B2(new_n223), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n239), .A2(KEYINPUT88), .A3(new_n240), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n245), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT93), .B1(new_n251), .B2(KEYINPUT17), .ZN(new_n252));
  OAI211_X1 g051(.A(KEYINPUT17), .B(new_n231), .C1(new_n237), .C2(new_n241), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n244), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n242), .A2(new_n218), .ZN(new_n257));
  NAND2_X1  g056(.A1(G229gat), .A2(G233gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(KEYINPUT18), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n218), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n251), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n257), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n258), .B(KEYINPUT13), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G197gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT11), .B(G169gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT12), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n254), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n249), .A2(new_n250), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n274), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(new_n231), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n259), .B1(new_n276), .B2(new_n244), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n272), .B1(new_n277), .B2(KEYINPUT18), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n202), .B1(new_n267), .B2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n277), .A2(KEYINPUT18), .B1(new_n264), .B2(new_n265), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT18), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n262), .B1(new_n251), .B2(KEYINPUT17), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n273), .B2(new_n275), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n283), .B2(new_n259), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(KEYINPUT94), .A3(new_n272), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n266), .A3(new_n261), .ZN(new_n287));
  INV_X1    g086(.A(new_n272), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT95), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n279), .A2(new_n285), .B1(new_n288), .B2(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT95), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G71gat), .B(G99gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT72), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(G15gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G43gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n303), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n307), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n311), .B1(new_n308), .B2(new_n309), .ZN(new_n312));
  OAI221_X1 g111(.A(new_n304), .B1(KEYINPUT28), .B2(new_n303), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n306), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n305), .B(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(KEYINPUT25), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(new_n302), .ZN(new_n323));
  AOI211_X1 g122(.A(new_n316), .B(new_n319), .C1(new_n320), .C2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n305), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n316), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n320), .A2(KEYINPUT65), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n320), .A2(KEYINPUT65), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n325), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n313), .B1(new_n324), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT1), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G113gat), .A2(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OR2_X1    g136(.A1(G127gat), .A2(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(G127gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT69), .B(G134gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G127gat), .B(G134gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n333), .A2(new_n334), .B1(KEYINPUT71), .B2(KEYINPUT1), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n342), .B(new_n343), .C1(KEYINPUT71), .C2(KEYINPUT1), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT70), .B(G120gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n332), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G227gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n348), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n300), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(KEYINPUT32), .C1(new_n355), .C2(new_n300), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n352), .B1(new_n349), .B2(new_n353), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT34), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI211_X1 g162(.A(KEYINPUT34), .B(new_n352), .C1(new_n349), .C2(new_n353), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n360), .A2(KEYINPUT73), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n360), .B2(KEYINPUT73), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(G22gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G141gat), .B(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(G155gat), .B2(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  XOR2_X1   g176(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G211gat), .B(G218gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT75), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT74), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n389), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n390));
  INV_X1    g189(.A(G197gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G204gat), .ZN(new_n392));
  INV_X1    g191(.A(G204gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G197gat), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n388), .A2(new_n390), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n383), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n383), .A2(new_n395), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT76), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n399), .A3(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n381), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n404), .A3(new_n400), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n377), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(G228gat), .B(G233gat), .C1(new_n403), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n375), .B(new_n376), .ZN(new_n410));
  INV_X1    g209(.A(new_n380), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n396), .B2(new_n397), .ZN(new_n412));
  INV_X1    g211(.A(new_n378), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n402), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n408), .B2(new_n415), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n371), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n422), .A2(new_n370), .A3(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n368), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n401), .ZN(new_n426));
  AND2_X1   g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n332), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n332), .A2(new_n404), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n426), .B(new_n428), .C1(new_n429), .C2(new_n427), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n427), .B1(new_n332), .B2(new_n380), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n401), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G8gat), .B(G36gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT78), .ZN(new_n435));
  XOR2_X1   g234(.A(G64gat), .B(G92gat), .Z(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT30), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n430), .B2(new_n433), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(KEYINPUT79), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n430), .A2(new_n433), .A3(new_n445), .A4(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n377), .A2(new_n348), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n379), .B(new_n347), .C1(new_n406), .C2(new_n377), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  XOR2_X1   g253(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n457), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n410), .B(new_n347), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n455), .A2(new_n452), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n459), .A2(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G1gat), .B(G29gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT0), .ZN(new_n465));
  XNOR2_X1  g264(.A(G57gat), .B(G85gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n449), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(new_n468), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT84), .B(new_n449), .C1(new_n463), .C2(new_n468), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n448), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n425), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  INV_X1    g277(.A(new_n472), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n475), .B1(new_n479), .B2(new_n469), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n360), .A2(new_n365), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n358), .B(new_n359), .C1(new_n363), .C2(new_n364), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n424), .ZN(new_n485));
  INV_X1    g284(.A(new_n448), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n477), .A2(new_n478), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n451), .A2(new_n453), .ZN(new_n490));
  INV_X1    g289(.A(new_n452), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n467), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n461), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT39), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n490), .B2(new_n491), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n489), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n472), .A2(new_n498), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n494), .A2(new_n497), .A3(new_n489), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n448), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n430), .A2(new_n433), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n438), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n428), .B1(new_n429), .B2(new_n427), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n401), .ZN(new_n506));
  OR3_X1    g305(.A1(new_n431), .A2(new_n432), .A3(new_n401), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT37), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT38), .ZN(new_n512));
  INV_X1    g311(.A(new_n502), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n511), .A2(new_n512), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n444), .A2(new_n446), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n516), .B(new_n475), .C1(new_n479), .C2(new_n469), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n501), .B(new_n485), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT36), .B1(new_n481), .B2(new_n482), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n368), .B2(KEYINPUT36), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n476), .A2(new_n485), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n296), .B1(new_n488), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(G57gat), .B2(G64gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G71gat), .A2(G78gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G71gat), .A2(G78gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT96), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G57gat), .ZN(new_n533));
  INV_X1    g332(.A(G64gat), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n528), .A2(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(G57gat), .A3(G64gat), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G57gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(KEYINPUT96), .ZN(new_n543));
  AND2_X1   g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n543), .A2(G64gat), .B1(new_n544), .B2(new_n527), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n538), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT97), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n531), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(new_n339), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n339), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n218), .B1(KEYINPUT21), .B2(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n556), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n556), .B2(new_n558), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G190gat), .B(G218gat), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT7), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(KEYINPUT98), .A3(G85gat), .A4(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578));
  NAND2_X1  g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(KEYINPUT8), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n576), .A2(new_n580), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT8), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(G99gat), .B2(G106gat), .ZN(new_n590));
  AND2_X1   g389(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n593), .B2(new_n582), .ZN(new_n594));
  INV_X1    g393(.A(new_n587), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n576), .A4(new_n580), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n242), .B2(new_n243), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n276), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n600));
  INV_X1    g399(.A(new_n597), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n251), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n571), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n571), .A3(new_n603), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n569), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g406(.A(new_n570), .B(new_n602), .C1(new_n276), .C2(new_n598), .ZN(new_n608));
  INV_X1    g407(.A(new_n569), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n565), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n531), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n540), .B1(new_n535), .B2(new_n539), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT97), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n588), .A3(new_n596), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n597), .A2(new_n548), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n548), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(KEYINPUT101), .A3(new_n622), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n618), .A2(new_n620), .ZN(new_n630));
  INV_X1    g429(.A(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n629), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n631), .B1(new_n621), .B2(new_n622), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n630), .B2(new_n631), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n638), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n613), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n524), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n474), .A2(new_n475), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n207), .ZN(G1324gat));
  OR3_X1    g444(.A1(new_n642), .A2(KEYINPUT102), .A3(new_n486), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT102), .B1(new_n642), .B2(new_n486), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(G8gat), .A3(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  NAND4_X1  g449(.A1(new_n649), .A2(KEYINPUT42), .A3(new_n448), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n646), .B2(new_n647), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n648), .B(new_n651), .C1(new_n653), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n642), .B2(new_n520), .ZN(new_n655));
  INV_X1    g454(.A(new_n483), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n655), .B1(new_n642), .B2(new_n657), .ZN(G1326gat));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n485), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT43), .B(G22gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  AOI21_X1  g460(.A(new_n478), .B1(new_n425), .B2(new_n476), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n487), .A2(new_n484), .ZN(new_n663));
  OAI22_X1  g462(.A1(new_n662), .A2(new_n663), .B1(new_n521), .B2(new_n522), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n611), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(KEYINPUT44), .A3(new_n611), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n565), .A2(new_n640), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n292), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G29gat), .B1(new_n673), .B2(new_n643), .ZN(new_n674));
  AND4_X1   g473(.A1(new_n664), .A2(new_n295), .A3(new_n611), .A4(new_n670), .ZN(new_n675));
  INV_X1    g474(.A(new_n643), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n224), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n225), .A3(new_n448), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT46), .Z(new_n681));
  OAI21_X1  g480(.A(G36gat), .B1(new_n673), .B2(new_n486), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(G1329gat));
  INV_X1    g482(.A(new_n520), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n667), .A2(new_n684), .A3(new_n668), .A4(new_n672), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n656), .A2(G43gat), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n675), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1330gat));
  NAND4_X1  g491(.A1(new_n667), .A2(new_n424), .A3(new_n668), .A4(new_n672), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g495(.A(G50gat), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n697), .A3(new_n424), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT48), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n693), .A2(G50gat), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n699), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n698), .A2(new_n700), .B1(KEYINPUT48), .B2(new_n702), .ZN(G1331gat));
  INV_X1    g502(.A(new_n613), .ZN(new_n704));
  AND4_X1   g503(.A1(new_n664), .A2(new_n292), .A3(new_n704), .A4(new_n640), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n643), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  INV_X1    g508(.A(KEYINPUT49), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n705), .B(new_n448), .C1(new_n710), .C2(new_n534), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n534), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  NAND2_X1  g512(.A1(new_n705), .A2(new_n684), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n656), .A2(G71gat), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n714), .A2(G71gat), .B1(new_n705), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n705), .A2(new_n424), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n565), .A2(new_n290), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n640), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n669), .A2(new_n676), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n612), .B1(new_n488), .B2(new_n523), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT51), .A4(new_n720), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n664), .A2(KEYINPUT51), .A3(new_n611), .A4(new_n720), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n665), .B2(new_n721), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n676), .A2(new_n593), .A3(new_n640), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n724), .A2(new_n593), .B1(new_n733), .B2(new_n734), .ZN(G1336gat));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n728), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n486), .A2(G92gat), .A3(new_n722), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n667), .A2(new_n448), .A3(new_n668), .A4(new_n723), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(G92gat), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT52), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n732), .A2(new_n737), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(new_n739), .B2(G92gat), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT107), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT107), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(G1337gat));
  NOR3_X1   g545(.A1(new_n656), .A2(G99gat), .A3(new_n722), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n667), .A2(new_n684), .A3(new_n668), .A4(new_n723), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G99gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(KEYINPUT108), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1338gat));
  NOR3_X1   g554(.A1(new_n485), .A2(G106gat), .A3(new_n722), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n732), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n667), .A2(new_n424), .A3(new_n668), .A4(new_n723), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G106gat), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n736), .A2(new_n756), .B1(new_n758), .B2(G106gat), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n757), .A2(new_n761), .B1(new_n762), .B2(new_n760), .ZN(G1339gat));
  NOR3_X1   g562(.A1(new_n613), .A2(new_n290), .A3(new_n640), .ZN(new_n764));
  INV_X1    g563(.A(new_n271), .ZN(new_n765));
  INV_X1    g564(.A(new_n265), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n263), .A2(new_n257), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n258), .ZN(new_n770));
  INV_X1    g569(.A(new_n257), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n283), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n765), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n286), .A2(new_n640), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n635), .B1(new_n637), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n621), .A2(new_n631), .A3(new_n622), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n631), .B1(new_n623), .B2(new_n624), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n627), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n778), .B1(new_n782), .B2(KEYINPUT109), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n784), .B(new_n780), .C1(new_n627), .C2(new_n781), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n776), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n628), .B2(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(KEYINPUT109), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n788), .A4(new_n778), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n636), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n775), .B1(new_n790), .B2(new_n292), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n612), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n611), .A2(new_n786), .A3(new_n636), .A4(new_n789), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n286), .A2(new_n774), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n286), .A2(KEYINPUT111), .A3(new_n774), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n563), .A2(new_n564), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n764), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n424), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n676), .A2(new_n486), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n656), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n333), .A3(new_n296), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n704), .A2(new_n292), .A3(new_n722), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT111), .B1(new_n286), .B2(new_n774), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n795), .B(new_n773), .C1(new_n279), .C2(new_n285), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n810), .A2(new_n793), .B1(new_n791), .B2(new_n612), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n565), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n707), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n368), .A2(new_n448), .A3(new_n424), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n290), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n806), .B1(new_n818), .B2(new_n333), .ZN(G1340gat));
  OAI21_X1  g618(.A(G120gat), .B1(new_n805), .B2(new_n722), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n640), .A2(new_n345), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT112), .Z(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n816), .B2(new_n822), .ZN(G1341gat));
  OAI21_X1  g622(.A(G127gat), .B1(new_n805), .B2(new_n800), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n565), .A2(new_n339), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n816), .B2(new_n825), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n817), .A2(new_n827), .A3(new_n340), .A4(new_n611), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n817), .A2(new_n340), .A3(new_n611), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n802), .A2(new_n611), .A3(new_n804), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n830), .A2(KEYINPUT56), .B1(new_n831), .B2(G134gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(G1343gat));
  NOR2_X1   g632(.A1(new_n803), .A2(new_n684), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n424), .A2(KEYINPUT57), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n786), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT114), .B(new_n776), .C1(new_n783), .C2(new_n785), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n789), .A2(new_n636), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI221_X4 g640(.A(KEYINPUT95), .B1(new_n288), .B2(new_n287), .C1(new_n279), .C2(new_n285), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n293), .B1(new_n286), .B2(new_n289), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n839), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n611), .B1(new_n844), .B2(new_n775), .ZN(new_n845));
  INV_X1    g644(.A(new_n798), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n800), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n835), .B1(new_n847), .B2(new_n807), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n812), .B2(new_n424), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n295), .B(new_n834), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n801), .B2(new_n485), .ZN(new_n853));
  INV_X1    g652(.A(new_n775), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n840), .B1(new_n837), .B2(new_n838), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n295), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n798), .B1(new_n856), .B2(new_n611), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n764), .B1(new_n857), .B2(new_n800), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n858), .B2(new_n835), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n295), .A4(new_n834), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n851), .A2(G141gat), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n813), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n812), .A2(KEYINPUT115), .A3(new_n707), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n684), .A2(new_n448), .A3(new_n485), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n296), .A2(G141gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n290), .B(new_n834), .C1(new_n848), .C2(new_n849), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G141gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n868), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(G141gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n850), .B2(KEYINPUT116), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n870), .B1(new_n880), .B2(new_n861), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n869), .B1(new_n875), .B2(new_n868), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT117), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n878), .A2(new_n883), .ZN(G1344gat));
  AND2_X1   g683(.A1(new_n864), .A2(new_n866), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n865), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n640), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n859), .A2(new_n640), .A3(new_n834), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n889), .A2(new_n890), .A3(G148gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n424), .A2(new_n852), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n641), .A2(new_n296), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n847), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n852), .B1(new_n812), .B2(new_n424), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n640), .A3(new_n834), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n888), .B1(new_n891), .B2(new_n898), .ZN(G1345gat));
  NAND4_X1  g698(.A1(new_n859), .A2(G155gat), .A3(new_n565), .A4(new_n834), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n565), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n885), .A2(KEYINPUT118), .A3(new_n565), .A4(new_n865), .ZN(new_n905));
  INV_X1    g704(.A(G155gat), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n904), .B2(new_n907), .ZN(G1346gat));
  INV_X1    g707(.A(G162gat), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n885), .A2(new_n909), .A3(new_n611), .A4(new_n865), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT119), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n859), .A2(new_n611), .A3(new_n834), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n801), .A2(new_n676), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n368), .A2(new_n486), .A3(new_n424), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(G169gat), .A3(new_n292), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT121), .Z(new_n921));
  NOR3_X1   g720(.A1(new_n707), .A2(new_n486), .A3(new_n656), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n802), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n296), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(G1348gat));
  OAI21_X1  g724(.A(G176gat), .B1(new_n923), .B2(new_n722), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n722), .A2(G176gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n919), .B2(new_n927), .ZN(G1349gat));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n565), .A2(new_n301), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n919), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n802), .A2(new_n922), .A3(new_n565), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n933), .A2(KEYINPUT122), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n322), .B1(new_n933), .B2(KEYINPUT122), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n923), .B2(new_n612), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n611), .A2(new_n302), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n919), .B2(new_n941), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n707), .A2(new_n486), .A3(new_n684), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n896), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n391), .A3(new_n296), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n520), .A2(new_n448), .A3(new_n424), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n917), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n290), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n945), .B1(new_n951), .B2(new_n391), .ZN(G1352gat));
  OAI21_X1  g751(.A(G204gat), .B1(new_n944), .B2(new_n722), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n640), .A2(new_n393), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT62), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n949), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n953), .A2(KEYINPUT126), .A3(new_n955), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1353gat));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n949), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n565), .A2(new_n385), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT127), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n966), .A3(new_n385), .A4(new_n565), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G211gat), .B1(new_n944), .B2(new_n800), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n944), .B2(new_n612), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n611), .A2(new_n386), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n963), .B2(new_n974), .ZN(G1355gat));
endmodule


