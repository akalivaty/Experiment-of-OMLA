//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND4_X1   g006(.A1(G143), .A2(new_n191), .A3(G214), .A4(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(G953), .B1(new_n188), .B2(new_n190), .ZN(new_n194));
  AOI21_X1  g008(.A(G143), .B1(new_n194), .B2(G214), .ZN(new_n195));
  OAI211_X1 g009(.A(KEYINPUT17), .B(G131), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT91), .ZN(new_n197));
  OAI21_X1  g011(.A(G131), .B1(new_n193), .B2(new_n195), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(G214), .A3(new_n192), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(G143), .A3(G214), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n199), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT16), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n212), .A3(G146), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n213), .B2(new_n214), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n204), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT17), .A4(G131), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n197), .A2(new_n206), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G113), .B(G122), .ZN(new_n223));
  INV_X1    g037(.A(G104), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n193), .A2(new_n195), .B1(new_n226), .B2(new_n203), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n203), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n202), .A2(new_n204), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT65), .B(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(G125), .B(G140), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n232), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT90), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n237));
  INV_X1    g051(.A(new_n235), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n237), .B(new_n238), .C1(new_n227), .C2(new_n229), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n222), .B(new_n225), .C1(new_n236), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n202), .A2(new_n204), .A3(new_n228), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n228), .B1(new_n202), .B2(new_n204), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n237), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n230), .A2(KEYINPUT90), .A3(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(KEYINPUT92), .A3(new_n225), .A4(new_n222), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n225), .B1(new_n248), .B2(new_n222), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n254));
  INV_X1    g068(.A(G902), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n242), .B2(new_n249), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT93), .B1(new_n257), .B2(G902), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(G475), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n198), .A2(new_n205), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n216), .B(KEYINPUT76), .Z(new_n261));
  INV_X1    g075(.A(new_n231), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n232), .B(KEYINPUT19), .Z(new_n263));
  OAI211_X1 g077(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n225), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n250), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n269));
  NOR2_X1   g083(.A1(G475), .A2(G902), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n242), .A2(new_n249), .B1(new_n266), .B2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(new_n270), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT20), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n259), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT94), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT94), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n259), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  XOR2_X1   g093(.A(G116), .B(G122), .Z(new_n280));
  OR2_X1    g094(.A1(KEYINPUT79), .A2(G107), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT79), .A2(G107), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT14), .A3(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G107), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G143), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT95), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT67), .B(G134), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n289), .A2(G143), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n291), .B2(new_n294), .ZN(new_n297));
  OAI221_X1 g111(.A(new_n284), .B1(new_n285), .B2(new_n288), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n301), .A2(KEYINPUT96), .B1(KEYINPUT13), .B2(new_n293), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n300), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT96), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n280), .A2(new_n283), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n295), .A2(new_n307), .B1(new_n284), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n307), .B2(new_n295), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n298), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G217), .A3(new_n192), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n311), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(G902), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT98), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT15), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G478), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n317), .A2(KEYINPUT98), .A3(new_n319), .A4(G478), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n317), .A2(KEYINPUT98), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G952), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(KEYINPUT99), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(KEYINPUT99), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n192), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(G234), .B2(G237), .ZN(new_n330));
  AOI211_X1 g144(.A(new_n192), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT21), .B(G898), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n277), .A2(new_n279), .A3(new_n325), .A4(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  INV_X1    g152(.A(G107), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(G104), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(KEYINPUT3), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n281), .A3(new_n282), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n338), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n201), .A2(G146), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n231), .B2(G143), .ZN(new_n351));
  AND2_X1   g165(.A1(KEYINPUT0), .A2(G128), .ZN(new_n352));
  NOR2_X1   g166(.A1(KEYINPUT0), .A2(G128), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n231), .A2(G143), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n201), .A2(G146), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n352), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(KEYINPUT80), .A2(G101), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT80), .A2(G101), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(new_n340), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n344), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n342), .A2(KEYINPUT81), .A3(new_n344), .A4(new_n363), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n345), .A2(new_n346), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(KEYINPUT82), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT82), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n360), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT11), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n292), .B2(G137), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n292), .A2(G137), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT68), .B(G137), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n375), .A2(new_n299), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G131), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(new_n203), .A3(new_n377), .A4(new_n380), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT1), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n356), .A2(new_n386), .A3(G128), .A4(new_n357), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n356), .A2(new_n357), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n289), .B1(new_n350), .B2(KEYINPUT1), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n283), .A2(new_n224), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n341), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n370), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT10), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n386), .B1(new_n231), .B2(G143), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n351), .B1(new_n396), .B2(new_n289), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n395), .B1(new_n397), .B2(new_n387), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n368), .A2(new_n369), .B1(G101), .B2(new_n392), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n394), .A2(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n374), .A2(new_n385), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G140), .ZN(new_n402));
  INV_X1    g216(.A(G227), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n385), .B1(new_n374), .B2(new_n400), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n374), .A2(new_n385), .A3(new_n400), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n390), .A2(new_n370), .A3(new_n393), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n397), .A2(new_n387), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n370), .B2(new_n393), .ZN(new_n412));
  OAI211_X1 g226(.A(KEYINPUT12), .B(new_n384), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n394), .B1(new_n411), .B2(new_n399), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT12), .B1(new_n415), .B2(new_n384), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n406), .A2(new_n408), .B1(new_n417), .B2(new_n405), .ZN(new_n418));
  OAI21_X1  g232(.A(G469), .B1(new_n418), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n316), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n405), .B1(new_n401), .B2(new_n407), .ZN(new_n421));
  INV_X1    g235(.A(new_n405), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n409), .B(new_n422), .C1(new_n414), .C2(new_n416), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(G469), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n337), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n397), .A2(new_n209), .A3(new_n387), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT86), .B1(new_n359), .B2(G125), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n433), .B(new_n209), .C1(new_n355), .C2(new_n358), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT87), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n431), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n430), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n441), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n430), .C1(new_n436), .C2(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G110), .B(G122), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT70), .B(G119), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G116), .ZN(new_n449));
  INV_X1    g263(.A(G119), .ZN(new_n450));
  OR3_X1    g264(.A1(new_n450), .A2(KEYINPUT71), .A3(G116), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT71), .B1(new_n450), .B2(G116), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT2), .B(G113), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n449), .A2(new_n454), .A3(new_n451), .A4(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n347), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n370), .A2(new_n371), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n370), .A2(KEYINPUT82), .A3(new_n371), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n370), .A2(new_n393), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n449), .A2(KEYINPUT5), .A3(new_n451), .A4(new_n452), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G113), .B1(new_n449), .B2(KEYINPUT5), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n447), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n459), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n372), .B2(new_n373), .ZN(new_n473));
  INV_X1    g287(.A(new_n470), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n446), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n446), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(KEYINPUT85), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT85), .B1(new_n477), .B2(new_n478), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n445), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n444), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n475), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n432), .A2(new_n435), .A3(new_n430), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n441), .A2(new_n482), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n468), .B1(new_n466), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n487), .B2(new_n466), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n465), .B1(new_n489), .B2(new_n457), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n446), .B(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(new_n469), .B2(new_n399), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n485), .A2(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n484), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n483), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n481), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n481), .B2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n429), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n335), .A2(new_n428), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n448), .B2(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n450), .A2(new_n289), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n448), .B2(new_n289), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n506), .B2(new_n503), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  OAI22_X1  g322(.A1(new_n507), .A2(G110), .B1(new_n508), .B2(new_n506), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n261), .A2(new_n509), .A3(new_n233), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n507), .A2(G110), .B1(new_n508), .B2(new_n506), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n215), .B2(new_n217), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT22), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(G137), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT77), .Z(new_n517));
  OR2_X1    g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G234), .ZN(new_n521));
  OAI21_X1  g335(.A(G217), .B1(new_n420), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n255), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n316), .A3(new_n519), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n525), .A2(KEYINPUT25), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n522), .B1(new_n525), .B2(KEYINPUT25), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n359), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n384), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n378), .A2(G134), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n292), .A2(G137), .ZN(new_n533));
  OAI21_X1  g347(.A(G131), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n383), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n411), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n536), .A3(KEYINPUT30), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(KEYINPUT69), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n383), .A2(new_n534), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n397), .B2(new_n387), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n382), .A2(new_n383), .B1(new_n359), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n530), .A2(KEYINPUT66), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n538), .A2(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n458), .B(new_n537), .C1(new_n545), .C2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n458), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n531), .A2(new_n536), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n194), .A2(G210), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT27), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT26), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n555), .A2(new_n556), .A3(G101), .ZN(new_n557));
  AOI21_X1  g371(.A(G101), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n548), .A2(new_n550), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n338), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n556), .A3(G101), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n550), .B(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n545), .A2(new_n549), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n548), .A2(new_n570), .A3(new_n559), .A4(new_n550), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n561), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n565), .A2(new_n550), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n548), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n559), .B1(new_n567), .B2(new_n568), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT29), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n549), .B1(new_n531), .B2(new_n536), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n567), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n559), .A2(KEYINPUT29), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n316), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n577), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n576), .A2(new_n586), .A3(KEYINPUT74), .A4(new_n577), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n529), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n502), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n363), .ZN(G3));
  NAND2_X1  g410(.A1(new_n427), .A2(new_n528), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n429), .B(new_n334), .C1(new_n498), .C2(new_n499), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n572), .A2(new_n316), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n574), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n315), .B(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G478), .A3(new_n316), .ZN(new_n604));
  INV_X1    g418(.A(G478), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n317), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n279), .B2(new_n277), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NOR2_X1   g426(.A1(new_n325), .A2(new_n276), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n335), .A2(new_n500), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n526), .A2(new_n527), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n517), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n513), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n255), .A3(new_n522), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n427), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n601), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n617), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT37), .B(G110), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G12));
  NAND2_X1  g442(.A1(new_n481), .A2(new_n496), .ZN(new_n629));
  INV_X1    g443(.A(new_n497), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n481), .A2(new_n496), .A3(new_n497), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(new_n427), .A3(new_n429), .A4(new_n623), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n589), .B2(new_n590), .ZN(new_n635));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n331), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n330), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n324), .A2(new_n259), .A3(new_n275), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  XNOR2_X1  g457(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT101), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n633), .B(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n429), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n623), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n259), .A2(new_n278), .A3(new_n275), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n278), .B1(new_n259), .B2(new_n275), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n325), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n576), .A2(new_n577), .ZN(new_n653));
  INV_X1    g467(.A(new_n578), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n255), .B1(new_n654), .B2(new_n582), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n565), .B1(new_n548), .B2(new_n550), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n648), .A2(new_n661), .A3(new_n652), .A4(new_n658), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n639), .B(KEYINPUT103), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT39), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n427), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT40), .Z(new_n666));
  AND3_X1   g480(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n201), .ZN(G45));
  OAI211_X1 g482(.A(new_n607), .B(new_n639), .C1(new_n649), .C2(new_n650), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n277), .A2(new_n279), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n607), .A4(new_n639), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n635), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT105), .B(G146), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G48));
  INV_X1    g490(.A(new_n598), .ZN(new_n677));
  INV_X1    g491(.A(new_n424), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(G469), .ZN(new_n680));
  INV_X1    g494(.A(G469), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT106), .B1(new_n424), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n336), .A3(new_n426), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n591), .A2(new_n609), .A3(new_n677), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT107), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n686), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n591), .A2(new_n677), .A3(new_n613), .A4(new_n685), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT108), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n286), .ZN(G18));
  INV_X1    g506(.A(new_n623), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n684), .A2(new_n500), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n589), .A2(new_n590), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n325), .A2(new_n334), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n649), .A3(new_n650), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  AOI21_X1  g513(.A(new_n647), .B1(new_n631), .B2(new_n632), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n324), .C1(new_n649), .C2(new_n650), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n583), .A2(new_n565), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n561), .A3(new_n571), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n573), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n600), .A2(new_n528), .A3(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n684), .A2(new_n706), .A3(new_n333), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  AND2_X1   g523(.A1(new_n600), .A2(new_n705), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n670), .A2(new_n673), .A3(new_n694), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n670), .A2(new_n673), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n427), .A2(new_n429), .A3(new_n631), .A4(new_n632), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n529), .B(new_n715), .C1(new_n589), .C2(new_n590), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n587), .A2(new_n528), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n715), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n670), .A2(new_n673), .A3(new_n718), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n714), .A2(new_n716), .B1(new_n719), .B2(KEYINPUT42), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  XNOR2_X1  g535(.A(new_n640), .B(KEYINPUT109), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NOR2_X1   g538(.A1(new_n633), .A2(new_n647), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n601), .A2(new_n623), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n671), .B(KEYINPUT110), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT43), .A3(new_n607), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n671), .B2(new_n608), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n725), .B1(new_n731), .B2(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(KEYINPUT44), .B2(new_n731), .ZN(new_n733));
  INV_X1    g547(.A(new_n426), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n418), .A2(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n418), .A2(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(G469), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(G469), .A2(G902), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n740), .B2(new_n739), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n336), .A3(new_n664), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n733), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT111), .B(G137), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G39));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n742), .A2(new_n747), .A3(new_n336), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n742), .B2(new_n336), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n725), .A2(new_n529), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n748), .A2(new_n749), .A3(new_n695), .A4(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n670), .A2(new_n673), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n207), .ZN(G42));
  NOR3_X1   g568(.A1(new_n608), .A2(new_n337), .A3(new_n647), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n734), .B1(new_n680), .B2(new_n682), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n755), .B(new_n528), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  INV_X1    g573(.A(new_n658), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n646), .A4(new_n727), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n649), .A2(new_n650), .A3(new_n325), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n602), .B1(new_n609), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n708), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n700), .A2(new_n757), .A3(new_n336), .A4(new_n623), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n335), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n695), .A2(new_n767), .B1(new_n617), .B2(new_n625), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n768), .A3(new_n686), .A4(new_n690), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n595), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n716), .A2(new_n713), .A3(new_n673), .A4(new_n670), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n723), .ZN(new_n773));
  INV_X1    g587(.A(new_n624), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n725), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n670), .A2(new_n673), .A3(new_n710), .ZN(new_n776));
  INV_X1    g590(.A(new_n639), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n276), .A2(new_n324), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n695), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n770), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n428), .A2(new_n623), .A3(new_n777), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n702), .A2(new_n658), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n711), .A2(new_n674), .A3(new_n642), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT52), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n762), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n674), .A2(new_n642), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n784), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n781), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n787), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n780), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n720), .A3(new_n723), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n626), .A2(new_n698), .A3(new_n764), .A4(new_n708), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n591), .A2(KEYINPUT78), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n501), .B1(new_n801), .B2(new_n592), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n802), .A3(new_n686), .A4(new_n690), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(KEYINPUT112), .A3(KEYINPUT53), .A4(new_n793), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n797), .A2(new_n787), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n795), .B1(KEYINPUT54), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n638), .B(new_n706), .C1(new_n728), .C2(new_n730), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n685), .A2(KEYINPUT113), .A3(new_n647), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT113), .B1(new_n685), .B2(new_n647), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n646), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n809), .A2(new_n813), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n638), .B1(new_n728), .B2(new_n730), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n757), .A2(new_n337), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n748), .B2(new_n749), .ZN(new_n822));
  INV_X1    g636(.A(new_n706), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n725), .ZN(new_n824));
  INV_X1    g638(.A(new_n725), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n684), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n623), .A3(new_n710), .A4(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n528), .A2(new_n826), .A3(new_n330), .A4(new_n760), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n651), .A3(new_n608), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n824), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n808), .B1(new_n819), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n329), .B1(new_n828), .B2(new_n609), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n820), .A2(new_n823), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n684), .A2(new_n500), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT116), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n832), .C1(new_n833), .C2(new_n835), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n820), .A2(new_n587), .A3(new_n528), .A4(new_n826), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT48), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(KEYINPUT48), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n837), .A2(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n830), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT51), .A3(new_n816), .A4(new_n818), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n831), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n807), .A2(KEYINPUT117), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n326), .A2(new_n192), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT117), .B1(new_n807), .B2(new_n846), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n761), .B1(new_n849), .B2(new_n850), .ZN(G75));
  NOR2_X1   g665(.A1(new_n192), .A2(G952), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n316), .B1(new_n787), .B2(new_n794), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n854), .B2(new_n630), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(new_n445), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT55), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n858), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(G51));
  NAND3_X1  g677(.A1(new_n787), .A2(new_n788), .A3(new_n794), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n787), .A2(new_n866), .A3(new_n788), .A4(new_n794), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n787), .A2(new_n794), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n738), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n421), .A2(new_n423), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n854), .A2(G469), .A3(new_n736), .A4(new_n735), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n852), .B1(new_n875), .B2(new_n876), .ZN(G54));
  NAND3_X1  g691(.A1(new_n854), .A2(KEYINPUT58), .A3(G475), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n878), .A2(new_n272), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n272), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n880), .A3(new_n852), .ZN(G60));
  NAND2_X1  g695(.A1(G478), .A2(G902), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT59), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n806), .A2(KEYINPUT54), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n864), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT121), .B1(new_n885), .B2(new_n603), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  INV_X1    g701(.A(new_n603), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(new_n807), .C2(new_n883), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n883), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n852), .B1(new_n870), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n886), .A2(new_n889), .A3(new_n891), .ZN(G63));
  NAND2_X1  g706(.A1(G217), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT60), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n520), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n621), .B(KEYINPUT122), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n896), .B(new_n853), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(G66));
  OAI21_X1  g714(.A(G953), .B1(new_n332), .B2(new_n440), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n803), .B2(new_n192), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n856), .B1(G898), .B2(new_n192), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n903), .B(new_n904), .Z(G69));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n801), .A2(new_n592), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n609), .A2(new_n763), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n907), .A2(new_n665), .A3(new_n908), .A4(new_n825), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n753), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n909), .A2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n744), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n789), .A2(new_n711), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n667), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n916), .A3(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n537), .B1(new_n545), .B2(new_n547), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n263), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n403), .A2(new_n636), .A3(new_n192), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n701), .A2(new_n717), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n743), .B1(new_n733), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n753), .A2(new_n913), .A3(new_n773), .ZN(new_n924));
  AOI21_X1  g738(.A(G953), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n403), .A2(G900), .A3(G953), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g741(.A1(new_n917), .A2(new_n921), .B1(new_n925), .B2(new_n927), .ZN(G72));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n579), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n656), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n806), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT127), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n579), .B(KEYINPUT126), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n923), .A2(new_n770), .A3(new_n924), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n930), .B(KEYINPUT125), .Z(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n912), .A2(new_n916), .A3(new_n803), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n656), .B1(new_n939), .B2(new_n937), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n853), .A2(new_n934), .A3(new_n938), .A4(new_n940), .ZN(G57));
endmodule


