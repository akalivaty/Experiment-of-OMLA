//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n196), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT73), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n200), .A2(KEYINPUT3), .B1(new_n201), .B2(G104), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  OAI22_X1  g018(.A1(KEYINPUT73), .A2(new_n203), .B1(new_n204), .B2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT3), .A4(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n207), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n207), .B2(new_n208), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n206), .ZN(new_n212));
  AOI22_X1  g026(.A1(KEYINPUT73), .A2(new_n203), .B1(new_n204), .B2(G107), .ZN(new_n213));
  AND4_X1   g027(.A1(new_n210), .A2(new_n212), .A3(new_n208), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT74), .B1(new_n207), .B2(new_n208), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT3), .A4(G104), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n200), .A2(KEYINPUT3), .B1(new_n201), .B2(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G101), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n221), .A3(KEYINPUT4), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n199), .B(new_n209), .C1(new_n215), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n201), .A2(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n204), .A2(G107), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n212), .A2(new_n208), .A3(new_n213), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT75), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n207), .A2(new_n210), .A3(new_n208), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT5), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(G113), .C1(KEYINPUT5), .C2(new_n192), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n197), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n223), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT79), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n223), .A2(new_n237), .A3(new_n233), .A4(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n234), .B1(new_n223), .B2(new_n233), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(KEYINPUT80), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n241), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT80), .B1(new_n239), .B2(new_n242), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT1), .B1(new_n249), .B2(G146), .ZN(new_n252));
  OAI21_X1  g066(.A(G128), .B1(new_n252), .B2(KEYINPUT67), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G143), .B2(new_n247), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n248), .A3(new_n250), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G143), .B(G146), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(KEYINPUT68), .B(new_n251), .C1(new_n253), .C2(new_n257), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT0), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n266), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n261), .A3(KEYINPUT64), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(KEYINPUT0), .B2(G128), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n274), .A2(new_n276), .B1(KEYINPUT0), .B2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n277), .B2(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G224), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n281), .B(new_n283), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n245), .A2(new_n246), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n232), .A2(new_n197), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n230), .B2(KEYINPUT82), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n230), .A2(KEYINPUT82), .A3(new_n287), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n234), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n281), .A2(new_n286), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n280), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n271), .B2(KEYINPUT83), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(KEYINPUT83), .B2(new_n271), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(new_n286), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n297), .B2(new_n239), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n190), .B1(new_n285), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n239), .A2(new_n242), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n284), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n303), .A2(new_n244), .A3(new_n243), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n298), .A3(new_n189), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n188), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT86), .B(G475), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT71), .A2(G125), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(KEYINPUT71), .A2(G125), .A3(G140), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT16), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n279), .B2(G140), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(new_n247), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n247), .B1(new_n314), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n282), .A3(G214), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(new_n249), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(KEYINPUT17), .A3(G131), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(G131), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n321), .B(G143), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n319), .B(new_n323), .C1(new_n328), .C2(KEYINPUT17), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT18), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n325), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n312), .A2(new_n313), .ZN(new_n333));
  MUX2_X1   g147(.A(new_n332), .B(new_n333), .S(G146), .Z(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(KEYINPUT18), .A3(G131), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT85), .B(G104), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n337), .B1(new_n342), .B2(new_n341), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n309), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT19), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n247), .A3(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n328), .A2(new_n347), .A3(new_n348), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n336), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n354), .A2(KEYINPUT84), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n341), .B1(new_n354), .B2(KEYINPUT84), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n338), .A2(new_n341), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n360));
  NOR2_X1   g174(.A1(G475), .A2(G902), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n355), .A2(new_n356), .B1(new_n338), .B2(new_n341), .ZN(new_n363));
  INV_X1    g177(.A(new_n361), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n346), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G478), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT15), .ZN(new_n369));
  INV_X1    g183(.A(G122), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G116), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n193), .A2(G122), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(new_n201), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n249), .A2(G128), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n249), .A2(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G134), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n373), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G116), .B2(new_n370), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(KEYINPUT90), .B2(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT89), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n389), .B2(new_n201), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT13), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n374), .B1(new_n391), .B2(new_n376), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n249), .A2(KEYINPUT13), .A3(G128), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n379), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n371), .A2(new_n372), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n201), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n395), .A2(new_n397), .A3(KEYINPUT88), .A4(new_n380), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n396), .A2(new_n201), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n380), .B1(new_n400), .B2(new_n373), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(new_n394), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  INV_X1    g217(.A(G217), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(G953), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n390), .A2(new_n398), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n201), .B1(new_n386), .B2(new_n388), .ZN(new_n407));
  INV_X1    g221(.A(new_n381), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n398), .B(new_n402), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI211_X1 g228(.A(KEYINPUT91), .B(G902), .C1(new_n406), .C2(new_n411), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n369), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n369), .B2(new_n414), .ZN(new_n417));
  INV_X1    g231(.A(G902), .ZN(new_n418));
  AOI211_X1 g232(.A(new_n418), .B(new_n282), .C1(G234), .C2(G237), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(KEYINPUT92), .A2(G952), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT92), .A2(G952), .ZN(new_n423));
  AOI21_X1  g237(.A(G953), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G234), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(new_n320), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n367), .A2(new_n417), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n307), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT26), .B(G101), .Z(new_n431));
  NAND3_X1  g245(.A1(new_n320), .A2(new_n282), .A3(G210), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT11), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n379), .B2(G137), .ZN(new_n438));
  INV_X1    g252(.A(G137), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT11), .A3(G134), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n438), .B(new_n440), .C1(G134), .C2(new_n439), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G131), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n379), .B2(G137), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(KEYINPUT65), .A3(G134), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(G134), .C2(new_n439), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n442), .B1(G131), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n269), .A2(new_n268), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n255), .A2(new_n256), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(G128), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT68), .B1(new_n451), .B2(new_n251), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n199), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n441), .B(G131), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n278), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n453), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT28), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n436), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n456), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT30), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n453), .A2(new_n467), .A3(new_n456), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n457), .B1(new_n469), .B2(new_n199), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT31), .B1(new_n470), .B2(new_n436), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n453), .A2(new_n467), .A3(new_n456), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n467), .B1(new_n453), .B2(new_n456), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n199), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n474), .A2(KEYINPUT31), .A3(new_n460), .A4(new_n436), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n464), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(G472), .A2(G902), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n459), .A2(new_n462), .A3(new_n436), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n436), .B1(new_n474), .B2(new_n460), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n418), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n459), .B2(new_n462), .ZN(new_n486));
  INV_X1    g300(.A(new_n458), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n460), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT70), .B1(new_n488), .B2(KEYINPUT28), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n436), .A2(KEYINPUT29), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n486), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G472), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n474), .A2(new_n460), .A3(new_n436), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT31), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n463), .B1(new_n496), .B2(new_n475), .ZN(new_n497));
  INV_X1    g311(.A(new_n478), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n479), .A2(new_n492), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n404), .B1(G234), .B2(new_n418), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n261), .A2(G119), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n261), .A2(KEYINPUT23), .A3(G119), .ZN(new_n506));
  INV_X1    g320(.A(G110), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n191), .A2(G128), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n503), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT24), .B(G110), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n509), .A2(new_n512), .B1(new_n247), .B2(new_n332), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n347), .A2(new_n348), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n508), .A3(new_n506), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G110), .ZN(new_n516));
  OAI221_X1 g330(.A(new_n516), .B1(new_n510), .B2(new_n511), .C1(new_n317), .C2(new_n318), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n282), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n517), .A3(new_n521), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n418), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(KEYINPUT25), .A3(new_n418), .A4(new_n524), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n502), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n524), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n521), .B1(new_n514), .B2(new_n517), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n501), .A2(G902), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n500), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G469), .ZN(new_n539));
  INV_X1    g353(.A(new_n226), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n251), .B1(new_n255), .B2(new_n261), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT66), .B1(new_n266), .B2(new_n262), .ZN(new_n542));
  AND4_X1   g356(.A1(KEYINPUT66), .A2(new_n262), .A3(new_n248), .A4(new_n250), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n540), .B(new_n544), .C1(new_n211), .C2(new_n214), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n270), .B2(new_n230), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n455), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT76), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT12), .B1(new_n455), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n278), .B(new_n209), .C1(new_n215), .C2(new_n222), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n270), .A2(KEYINPUT10), .A3(new_n230), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n455), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n552), .A2(new_n553), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n282), .A2(G227), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n546), .A2(new_n455), .A3(new_n549), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n551), .A2(new_n557), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n455), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n563), .A2(new_n564), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n539), .B(new_n418), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n563), .A2(new_n564), .B1(new_n568), .B2(new_n560), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n549), .B1(new_n546), .B2(new_n455), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n552), .A2(new_n555), .A3(new_n553), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(new_n556), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(KEYINPUT77), .A3(new_n561), .A4(new_n562), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n539), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n560), .A3(new_n562), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n568), .A2(new_n561), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G469), .B1(new_n585), .B2(G902), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n538), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n430), .A2(new_n536), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT93), .B(G101), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G3));
  AND3_X1   g404(.A1(new_n305), .A2(new_n298), .A3(new_n189), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n189), .B1(new_n305), .B2(new_n298), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n406), .A2(new_n411), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n406), .A2(new_n411), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n368), .A2(new_n418), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n412), .B2(new_n368), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n367), .ZN(new_n604));
  NOR4_X1   g418(.A1(new_n593), .A2(new_n188), .A3(new_n428), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(KEYINPUT94), .A2(G472), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n477), .A2(new_n418), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n497), .B2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(new_n529), .A3(new_n534), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n587), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT95), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  XOR2_X1   g429(.A(new_n427), .B(KEYINPUT96), .Z(new_n616));
  NAND3_X1  g430(.A1(new_n417), .A2(new_n366), .A3(new_n616), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n188), .B(new_n617), .C1(new_n300), .C2(new_n306), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n587), .A3(new_n611), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n527), .A2(new_n528), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n501), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n518), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n533), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n622), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n627), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n529), .A2(new_n629), .A3(KEYINPUT97), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n607), .A2(new_n631), .A3(new_n609), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n430), .A2(new_n633), .A3(new_n587), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n419), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n426), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT99), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n417), .A2(new_n366), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n187), .C1(new_n591), .C2(new_n592), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT100), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n300), .A2(new_n306), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n187), .A4(new_n642), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n500), .A2(new_n631), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n647), .A3(new_n587), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XOR2_X1   g464(.A(new_n640), .B(KEYINPUT39), .Z(new_n651));
  NAND2_X1  g465(.A1(new_n587), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT40), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n652), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT101), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n593), .B(KEYINPUT38), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n470), .A2(new_n435), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n418), .B1(new_n488), .B2(new_n436), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n479), .A2(new_n499), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n367), .A2(new_n417), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n529), .A2(new_n629), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n187), .A3(new_n667), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n659), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n655), .A2(new_n658), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  NOR3_X1   g485(.A1(new_n602), .A2(new_n366), .A3(new_n640), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n587), .A2(new_n648), .A3(new_n307), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NAND3_X1  g488(.A1(new_n578), .A2(new_n569), .A3(new_n565), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n539), .B1(new_n675), .B2(new_n418), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n580), .B1(new_n579), .B2(new_n539), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n580), .A2(new_n675), .A3(new_n539), .A4(new_n418), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n537), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n500), .A2(new_n535), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n605), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT41), .B(G113), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT102), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n683), .B(new_n685), .ZN(G15));
  AOI21_X1  g500(.A(new_n676), .B1(new_n573), .B2(new_n581), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n500), .A3(new_n535), .A4(new_n537), .ZN(new_n688));
  INV_X1    g502(.A(new_n617), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n645), .A2(new_n187), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT103), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n692));
  AOI211_X1 g506(.A(new_n538), .B(new_n676), .C1(new_n573), .C2(new_n581), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n618), .A2(new_n692), .A3(new_n536), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND4_X1  g510(.A1(new_n687), .A2(new_n645), .A3(new_n537), .A4(new_n187), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n429), .A2(new_n500), .A3(new_n631), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n698), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n693), .A4(new_n307), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n535), .B(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n497), .B2(G902), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n435), .B1(new_n486), .B2(new_n489), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n471), .B2(new_n476), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n478), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n706), .A2(new_n616), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n680), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n593), .A2(new_n188), .A3(new_n665), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  INV_X1    g529(.A(new_n667), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n710), .A2(new_n707), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n693), .A2(new_n307), .A3(new_n672), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  NOR3_X1   g533(.A1(new_n591), .A2(new_n592), .A3(new_n188), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n587), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n500), .A2(new_n706), .ZN(new_n722));
  INV_X1    g536(.A(new_n672), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n587), .A2(new_n536), .A3(new_n672), .A4(new_n720), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n724), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n728), .A2(KEYINPUT106), .A3(new_n724), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n326), .ZN(G33));
  NAND4_X1  g548(.A1(new_n587), .A2(new_n536), .A3(new_n642), .A4(new_n720), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G134), .ZN(G36));
  NAND2_X1  g550(.A1(new_n610), .A2(new_n716), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT108), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n367), .A2(new_n602), .A3(KEYINPUT43), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n603), .B1(new_n740), .B2(new_n366), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n367), .A2(KEYINPUT107), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n739), .B1(new_n743), .B2(KEYINPUT43), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n738), .A2(new_n744), .A3(KEYINPUT44), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT44), .B1(new_n738), .B2(new_n744), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n585), .A2(KEYINPUT45), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n585), .A2(KEYINPUT45), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n748), .A3(new_n539), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n539), .A2(new_n418), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n582), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n537), .A3(new_n651), .A4(new_n720), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n745), .A2(new_n746), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n439), .ZN(G39));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n537), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(KEYINPUT47), .A3(new_n537), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n720), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n763), .A2(new_n723), .A3(new_n500), .A4(new_n535), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT109), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n767), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  AOI22_X1  g584(.A1(new_n605), .A2(new_n682), .B1(new_n712), .B2(new_n713), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n703), .A2(new_n695), .A3(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n430), .B(new_n587), .C1(new_n633), .C2(new_n536), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n417), .A2(new_n366), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n604), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(new_n616), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n587), .A3(new_n307), .A4(new_n611), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n717), .A2(new_n672), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n367), .A2(new_n417), .A3(new_n640), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n500), .A3(new_n631), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n587), .A3(new_n720), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n773), .A2(new_n735), .A3(new_n777), .A4(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n733), .A2(new_n772), .A3(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n663), .A2(new_n667), .A3(new_n641), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n713), .A2(new_n587), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n649), .A2(new_n786), .A3(new_n673), .A4(new_n718), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n649), .A2(new_n718), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n787), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n784), .A2(KEYINPUT53), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n772), .A2(new_n783), .ZN(new_n794));
  INV_X1    g608(.A(new_n732), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT106), .B1(new_n728), .B2(new_n724), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n726), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n790), .A2(new_n788), .A3(new_n673), .A4(new_n786), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n793), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n800), .B2(new_n791), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT111), .B1(new_n800), .B2(new_n801), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  INV_X1    g622(.A(new_n801), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n784), .A2(new_n808), .A3(new_n789), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n804), .B1(KEYINPUT54), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n426), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n744), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n693), .A2(new_n720), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n717), .ZN(new_n817));
  INV_X1    g631(.A(new_n815), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n818), .A2(new_n535), .A3(new_n813), .A4(new_n664), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n602), .A2(new_n366), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n817), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n687), .A2(new_n538), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n760), .A2(new_n761), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n814), .A2(new_n824), .A3(new_n763), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n659), .A2(new_n188), .A3(new_n693), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n814), .A2(new_n824), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT50), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n834));
  OAI211_X1 g648(.A(new_n826), .B(new_n833), .C1(new_n831), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n830), .A2(new_n307), .A3(new_n693), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n424), .C1(new_n819), .C2(new_n604), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n816), .A2(new_n500), .A3(new_n706), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(KEYINPUT48), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(KEYINPUT48), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT115), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n812), .A2(new_n837), .A3(new_n838), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(G952), .B2(G953), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n706), .A2(new_n537), .A3(new_n187), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n743), .A2(new_n663), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n687), .B(KEYINPUT49), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n659), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(G75));
  AOI21_X1  g667(.A(new_n418), .B1(new_n793), .B2(new_n802), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(G210), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n284), .B1(new_n245), .B2(new_n246), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n305), .ZN(new_n859));
  XNOR2_X1  g673(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n859), .B(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n857), .A2(new_n861), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n282), .A2(G952), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G51));
  NAND2_X1  g679(.A1(new_n793), .A2(new_n802), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(G902), .A3(new_n749), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n854), .A2(new_n869), .A3(new_n749), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n675), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n793), .A2(new_n802), .A3(new_n803), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n751), .B(KEYINPUT57), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n873), .B2(new_n874), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT117), .B1(new_n881), .B2(new_n872), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n864), .B1(new_n879), .B2(new_n882), .ZN(G54));
  AND2_X1   g697(.A1(KEYINPUT58), .A2(G475), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n854), .A2(new_n359), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n359), .B1(new_n854), .B2(new_n884), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n864), .ZN(G60));
  XNOR2_X1  g701(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n600), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n874), .ZN(new_n891));
  INV_X1    g705(.A(new_n598), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT120), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n598), .C1(new_n812), .C2(new_n889), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n598), .A2(new_n889), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n864), .B1(new_n875), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(G63));
  INV_X1    g712(.A(new_n864), .ZN(new_n899));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT60), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n866), .A2(new_n626), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n866), .A2(new_n901), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n899), .B(new_n902), .C1(new_n903), .C2(new_n532), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n904), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT61), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G66));
  INV_X1    g721(.A(G224), .ZN(new_n908));
  OAI21_X1  g722(.A(G953), .B1(new_n420), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n773), .A2(new_n777), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n772), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(G953), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n245), .A2(new_n246), .B1(G898), .B2(new_n282), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G69));
  NAND2_X1  g728(.A1(new_n349), .A2(new_n351), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n469), .B(new_n915), .Z(new_n916));
  NAND2_X1  g730(.A1(G900), .A2(G953), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n797), .A2(new_n735), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT125), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n790), .A2(new_n673), .ZN(new_n920));
  INV_X1    g734(.A(new_n713), .ZN(new_n921));
  INV_X1    g735(.A(new_n651), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n758), .A2(new_n921), .A3(new_n922), .A4(new_n722), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n756), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n769), .A3(new_n920), .A4(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n916), .B(new_n917), .C1(new_n925), .C2(G953), .ZN(new_n926));
  INV_X1    g740(.A(new_n756), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n536), .A2(new_n720), .A3(new_n775), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n652), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT122), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n930), .A3(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n929), .B(KEYINPUT122), .Z(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(new_n756), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n670), .A2(new_n920), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n670), .A2(new_n938), .A3(new_n920), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n937), .A3(new_n769), .A4(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n931), .A2(new_n934), .B1(new_n766), .B2(new_n768), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n939), .A4(new_n937), .ZN(new_n944));
  AOI21_X1  g758(.A(G953), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n926), .B1(new_n945), .B2(new_n916), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n282), .B1(G227), .B2(G900), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n926), .B(new_n949), .C1(new_n945), .C2(new_n916), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G72));
  NAND3_X1  g767(.A1(new_n942), .A2(new_n911), .A3(new_n944), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI211_X1 g770(.A(new_n435), .B(new_n470), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n911), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n925), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n435), .A3(new_n470), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n494), .A2(KEYINPUT127), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(new_n483), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n811), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n899), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n957), .A2(new_n964), .ZN(G57));
endmodule


