//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n199), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n200), .A2(new_n202), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n187), .B1(new_n198), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n195), .A2(new_n197), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(G146), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n208), .B1(new_n219), .B2(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n214), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n218), .A2(new_n221), .A3(KEYINPUT69), .A4(new_n207), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G134), .B(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n224), .B2(new_n196), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n189), .A2(G137), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n191), .A2(G134), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n226), .B(G131), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n197), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT70), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n225), .A2(new_n232), .A3(new_n229), .A4(new_n197), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n219), .B2(G143), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT67), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT67), .A2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n220), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n203), .A2(new_n205), .A3(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n231), .A2(new_n233), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT2), .A2(G113), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT68), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT2), .A3(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT2), .A2(G113), .ZN(new_n249));
  XNOR2_X1  g063(.A(G116), .B(G119), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n248), .B2(new_n249), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT71), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n249), .ZN(new_n256));
  INV_X1    g070(.A(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n223), .A2(new_n243), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT72), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n254), .A2(new_n259), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n231), .A2(new_n233), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n238), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n242), .B1(new_n271), .B2(new_n212), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n273), .A3(new_n217), .A4(new_n222), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n266), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n273), .A2(KEYINPUT30), .A3(new_n217), .A4(new_n222), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n216), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n221), .A2(KEYINPUT65), .A3(new_n207), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n198), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n272), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n230), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n278), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n252), .A2(new_n253), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n277), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n268), .A2(new_n276), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n268), .A2(KEYINPUT31), .A3(new_n276), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n282), .B2(new_n284), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n274), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT28), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  OAI22_X1  g111(.A1(new_n254), .A2(new_n259), .B1(new_n198), .B2(new_n216), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n243), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n266), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n300), .B1(new_n291), .B2(new_n292), .ZN(new_n307));
  INV_X1    g121(.A(new_n303), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n299), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n223), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n269), .B1(new_n312), .B2(new_n273), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT28), .B1(new_n313), .B2(new_n261), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT29), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n297), .B1(new_n274), .B2(new_n294), .ZN(new_n317));
  INV_X1    g131(.A(new_n299), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n267), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n288), .A2(new_n274), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n316), .A3(new_n267), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT75), .B(G902), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G472), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n304), .A2(new_n309), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n304), .A2(new_n309), .A3(KEYINPUT76), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G217), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n323), .B2(G234), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G902), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n240), .A2(G119), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n238), .B2(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  INV_X1    g154(.A(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(G125), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n342), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n199), .ZN(new_n348));
  OAI211_X1 g162(.A(G146), .B(new_n342), .C1(new_n346), .C2(new_n340), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT23), .B1(new_n240), .B2(G119), .ZN(new_n351));
  INV_X1    g165(.A(G119), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(G128), .ZN(new_n353));
  OR2_X1    g167(.A1(KEYINPUT67), .A2(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT67), .A2(G128), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n354), .A2(KEYINPUT23), .A3(G119), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G110), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(KEYINPUT78), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n339), .B(new_n350), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n346), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n219), .ZN(new_n363));
  INV_X1    g177(.A(G110), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n353), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n336), .A2(new_n338), .B1(new_n365), .B2(KEYINPUT79), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n349), .B(new_n363), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G137), .ZN(new_n369));
  INV_X1    g183(.A(G953), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n370), .A2(G221), .A3(G234), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n369), .B(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n361), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n361), .B2(new_n368), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT81), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n361), .A2(new_n368), .ZN(new_n377));
  INV_X1    g191(.A(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n361), .A2(new_n368), .A3(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n333), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT82), .B(new_n333), .C1(new_n375), .C2(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n386));
  NOR2_X1   g200(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n380), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(new_n323), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n323), .B(new_n387), .C1(new_n373), .C2(new_n374), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n386), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n384), .A2(new_n385), .B1(new_n392), .B2(new_n332), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT17), .B(G131), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n348), .A2(new_n397), .A3(new_n349), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n348), .A2(new_n397), .A3(KEYINPUT91), .A4(new_n349), .ZN(new_n401));
  OAI21_X1  g215(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n370), .A3(G214), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n211), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n196), .A3(new_n394), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n402), .A2(KEYINPUT92), .A3(new_n403), .A4(new_n407), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n400), .A2(new_n401), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G113), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n363), .B1(new_n199), .B2(new_n362), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n406), .B(new_n394), .C1(new_n417), .C2(new_n196), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n416), .B(new_n418), .C1(new_n417), .C2(new_n402), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n402), .A2(new_n407), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n346), .B(KEYINPUT19), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n349), .B1(new_n422), .B2(new_n210), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n415), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT20), .ZN(new_n431));
  INV_X1    g245(.A(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n420), .B2(new_n426), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT93), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND4_X1   g249(.A1(KEYINPUT94), .A2(new_n427), .A3(new_n434), .A4(new_n428), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT94), .B1(new_n433), .B2(new_n434), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n431), .B(new_n435), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n420), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n415), .B1(new_n412), .B2(new_n419), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G475), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n236), .A2(new_n237), .A3(new_n211), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n240), .A2(G143), .ZN(new_n446));
  OAI21_X1  g260(.A(G134), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n354), .A2(G143), .A3(new_n355), .ZN(new_n448));
  INV_X1    g262(.A(new_n446), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n189), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G107), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT95), .B1(new_n452), .B2(G116), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT95), .ZN(new_n454));
  INV_X1    g268(.A(G116), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G122), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n453), .A2(new_n456), .B1(G116), .B2(new_n452), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n447), .A2(new_n450), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n455), .B2(G122), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n452), .A2(KEYINPUT95), .A3(G116), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(G116), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT9), .B(G234), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n468), .A2(new_n331), .A3(G953), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT96), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n448), .A2(KEYINPUT13), .A3(new_n449), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n189), .B1(new_n446), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n453), .A2(new_n456), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n476), .A2(new_n451), .A3(new_n462), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n451), .B1(new_n476), .B2(new_n462), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n475), .B(new_n450), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n467), .A2(new_n471), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n471), .B1(new_n467), .B2(new_n479), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT98), .B(new_n323), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n483), .A2(KEYINPUT97), .ZN(new_n485));
  INV_X1    g299(.A(G478), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n465), .A2(G107), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n457), .A2(new_n451), .ZN(new_n490));
  INV_X1    g304(.A(new_n450), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n189), .B1(new_n448), .B2(new_n449), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n479), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n471), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n467), .A2(new_n471), .A3(new_n479), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT98), .B1(new_n498), .B2(new_n323), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  AOI211_X1 g314(.A(KEYINPUT98), .B(new_n487), .C1(new_n498), .C2(new_n323), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT99), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G952), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(G953), .ZN(new_n504));
  INV_X1    g318(.A(G234), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(new_n404), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n370), .B(new_n323), .C1(G234), .C2(G237), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT21), .B(G898), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n323), .B1(new_n480), .B2(new_n481), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT98), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n482), .A3(new_n487), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n488), .A2(new_n499), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n502), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n444), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G469), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT10), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n204), .B1(new_n219), .B2(G143), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n240), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n242), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT83), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT3), .B1(new_n414), .B2(G107), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT3), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n451), .A3(G104), .ZN(new_n529));
  INV_X1    g343(.A(G101), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n414), .A2(G107), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n451), .A2(G104), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n414), .A2(G107), .ZN(new_n534));
  OAI21_X1  g348(.A(G101), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n525), .A2(new_n526), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n526), .B1(new_n525), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n522), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G101), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT4), .A3(new_n532), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n544), .A3(G101), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n543), .A2(new_n207), .A3(new_n221), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n536), .A2(new_n522), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n272), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n540), .A2(new_n549), .A3(new_n198), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT84), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n540), .A2(new_n549), .A3(KEYINPUT84), .A4(new_n198), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI22_X1  g368(.A1(new_n538), .A2(new_n539), .B1(new_n272), .B2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n218), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G140), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n370), .A2(G227), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n561), .B(new_n562), .Z(new_n563));
  AND3_X1   g377(.A1(new_n554), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n540), .A2(new_n549), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n218), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n554), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n521), .B(new_n323), .C1(new_n564), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n554), .A2(new_n560), .ZN(new_n569));
  INV_X1    g383(.A(new_n563), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n570), .B1(new_n552), .B2(new_n553), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n566), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(G469), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n521), .A2(new_n439), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n568), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G221), .B1(new_n468), .B2(G902), .ZN(new_n578));
  OAI21_X1  g392(.A(G214), .B1(G237), .B2(G902), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n579), .B(KEYINPUT85), .Z(new_n580));
  OAI21_X1  g394(.A(G210), .B1(G237), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n583));
  XNOR2_X1  g397(.A(G110), .B(G122), .ZN(new_n584));
  XOR2_X1   g398(.A(new_n584), .B(KEYINPUT8), .Z(new_n585));
  INV_X1    g399(.A(KEYINPUT86), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n352), .A2(G116), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(KEYINPUT5), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n455), .A2(G119), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n589), .A3(KEYINPUT5), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT5), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n591), .A2(new_n352), .A3(KEYINPUT86), .A4(G116), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n588), .A2(new_n590), .A3(G113), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n251), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT88), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT88), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n596), .A3(new_n251), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n536), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n536), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT89), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n593), .A2(new_n596), .A3(new_n251), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n593), .B2(new_n251), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n537), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT89), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n585), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n370), .A2(G224), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT87), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT7), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n221), .A2(G125), .A3(new_n207), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(G125), .B1(new_n239), .B2(new_n242), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n272), .A2(new_n344), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n615), .A2(KEYINPUT7), .A3(new_n609), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n537), .A2(new_n251), .A3(new_n593), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n543), .A2(new_n545), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n584), .B(new_n618), .C1(new_n619), .C2(new_n286), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n583), .B(new_n439), .C1(new_n607), .C2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n618), .B1(new_n619), .B2(new_n286), .ZN(new_n623));
  INV_X1    g437(.A(new_n584), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n620), .A3(KEYINPUT6), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT6), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n623), .A2(new_n627), .A3(new_n624), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n629));
  INV_X1    g443(.A(new_n609), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n615), .A2(new_n630), .A3(new_n611), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n626), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n622), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n585), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n605), .B1(new_n604), .B2(new_n599), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n595), .A2(new_n597), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT89), .B1(new_n637), .B2(new_n537), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n623), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n584), .A2(new_n640), .B1(new_n614), .B2(new_n616), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n583), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n582), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n626), .A2(new_n628), .A3(new_n632), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n642), .B2(new_n583), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n439), .B1(new_n607), .B2(new_n621), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT90), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n646), .A2(new_n581), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n580), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n520), .A2(new_n577), .A3(new_n578), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n330), .A2(new_n393), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G101), .ZN(G3));
  INV_X1    g468(.A(new_n323), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n486), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT33), .B1(new_n480), .B2(new_n481), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT33), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n496), .A2(new_n659), .A3(new_n497), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(G478), .B1(new_n498), .B2(new_n323), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(KEYINPUT100), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n661), .B2(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n438), .B2(new_n443), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n650), .A3(new_n511), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n302), .A2(new_n303), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n307), .B2(new_n655), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n393), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n577), .A2(new_n578), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT34), .B(G104), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  XNOR2_X1  g491(.A(new_n443), .B(KEYINPUT101), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n431), .B(new_n435), .C1(KEYINPUT20), .C2(new_n429), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n502), .A2(new_n518), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n511), .A3(new_n650), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n577), .A2(new_n578), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n671), .A2(new_n672), .A3(new_n393), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NOR2_X1   g502(.A1(new_n372), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT102), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n377), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n333), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n373), .A2(new_n374), .ZN(new_n693));
  OAI22_X1  g507(.A1(new_n693), .A2(new_n655), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n694), .A2(new_n390), .B1(KEYINPUT80), .B2(KEYINPUT25), .ZN(new_n695));
  INV_X1    g509(.A(new_n332), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n671), .A2(new_n672), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n684), .A3(new_n520), .A4(new_n650), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(new_n508), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n506), .B1(new_n702), .B2(G900), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT103), .Z(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n650), .A2(new_n682), .A3(new_n697), .A4(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n674), .B1(new_n328), .B2(new_n329), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XOR2_X1   g523(.A(new_n704), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n684), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  INV_X1    g527(.A(new_n580), .ZN(new_n714));
  INV_X1    g528(.A(G472), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n267), .B1(new_n313), .B2(new_n261), .ZN(new_n716));
  AOI21_X1  g530(.A(G902), .B1(new_n289), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n304), .B(new_n309), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n697), .ZN(new_n719));
  INV_X1    g533(.A(new_n444), .ZN(new_n720));
  INV_X1    g534(.A(new_n681), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n714), .A2(new_n718), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n644), .A2(new_n649), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT38), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n712), .A2(new_n713), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NAND2_X1  g541(.A1(new_n669), .A2(new_n705), .ZN(new_n728));
  INV_X1    g542(.A(new_n650), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n728), .A2(new_n719), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n330), .A2(new_n684), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n707), .A2(new_n733), .A3(new_n730), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n554), .A2(new_n566), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n738), .A2(new_n570), .B1(new_n572), .B2(new_n560), .ZN(new_n739));
  OAI21_X1  g553(.A(G469), .B1(new_n739), .B2(new_n655), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n568), .ZN(new_n742));
  OAI211_X1 g556(.A(KEYINPUT105), .B(G469), .C1(new_n739), .C2(new_n655), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n737), .B1(new_n744), .B2(new_n578), .ZN(new_n745));
  INV_X1    g559(.A(new_n578), .ZN(new_n746));
  AOI211_X1 g560(.A(KEYINPUT106), .B(new_n746), .C1(new_n742), .C2(new_n743), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n393), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n328), .B2(new_n329), .ZN(new_n750));
  INV_X1    g564(.A(new_n670), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NAND3_X1  g568(.A1(new_n748), .A2(new_n683), .A3(new_n750), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT107), .B(G116), .Z(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G18));
  NAND2_X1  g571(.A1(new_n520), .A2(new_n697), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n328), .B2(new_n329), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n748), .A2(new_n650), .A3(new_n759), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT108), .B(G119), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G21));
  NAND3_X1  g576(.A1(new_n722), .A2(new_n511), .A3(new_n650), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n311), .A2(new_n314), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n293), .B1(new_n764), .B2(new_n266), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n303), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n393), .A3(new_n672), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n748), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G122), .ZN(G24));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n672), .A3(new_n697), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n728), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n748), .A2(new_n650), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  INV_X1    g588(.A(new_n728), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n644), .A2(new_n649), .A3(new_n714), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n574), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n569), .A2(new_n570), .B1(new_n572), .B2(new_n566), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT109), .A3(G469), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n568), .A2(new_n576), .ZN(new_n782));
  AOI211_X1 g596(.A(new_n746), .B(new_n776), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n330), .A2(new_n393), .A3(new_n775), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n784), .A2(KEYINPUT110), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT110), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n304), .A2(KEYINPUT111), .ZN(new_n788));
  INV_X1    g602(.A(new_n671), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n788), .B(new_n325), .C1(KEYINPUT32), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n304), .A2(KEYINPUT111), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n393), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n775), .ZN(new_n793));
  OAI22_X1  g607(.A1(new_n786), .A2(new_n787), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  NAND4_X1  g609(.A1(new_n750), .A2(new_n682), .A3(new_n705), .A4(new_n783), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g612(.A1(KEYINPUT45), .A2(G469), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n574), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT112), .B(G469), .C1(new_n779), .C2(KEYINPUT45), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n779), .A2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT46), .B(new_n576), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n805), .A2(new_n806), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n575), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n803), .B(new_n804), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(KEYINPUT114), .A3(KEYINPUT46), .A4(new_n576), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(new_n812), .A3(new_n814), .A4(new_n568), .ZN(new_n815));
  INV_X1    g629(.A(new_n776), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n444), .A2(KEYINPUT43), .A3(new_n668), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT43), .B1(new_n444), .B2(new_n668), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n671), .A2(new_n672), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n697), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n816), .B1(new_n822), .B2(KEYINPUT44), .ZN(new_n823));
  INV_X1    g637(.A(new_n819), .ZN(new_n824));
  INV_X1    g638(.A(new_n821), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n822), .A2(KEYINPUT115), .A3(KEYINPUT44), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n815), .A2(new_n830), .A3(new_n578), .A4(new_n710), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G137), .ZN(G39));
  NOR4_X1   g646(.A1(new_n330), .A2(new_n393), .A3(new_n728), .A4(new_n776), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT116), .Z(new_n834));
  NAND2_X1  g648(.A1(new_n815), .A2(new_n578), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT47), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n578), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(new_n341), .ZN(G42));
  NAND2_X1  g654(.A1(new_n824), .A2(new_n507), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n767), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n816), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT123), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n837), .A2(new_n838), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n578), .B1(new_n742), .B2(new_n743), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n745), .A2(new_n747), .A3(new_n776), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n718), .A2(new_n749), .A3(new_n506), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n720), .A3(new_n668), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n507), .A3(new_n824), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n841), .A2(new_n725), .A3(new_n714), .A4(new_n767), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n852), .A2(KEYINPUT50), .A3(new_n748), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT50), .B1(new_n852), .B2(new_n748), .ZN(new_n854));
  OAI221_X1 g668(.A(new_n850), .B1(new_n771), .B2(new_n851), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n847), .A2(KEYINPUT51), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n851), .A2(new_n792), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT48), .Z(new_n859));
  NAND3_X1  g673(.A1(new_n848), .A2(new_n669), .A3(new_n849), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n745), .A2(new_n747), .A3(new_n729), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n503), .B(G953), .C1(new_n842), .C2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n847), .B2(new_n856), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n794), .A2(new_n796), .ZN(new_n866));
  AOI211_X1 g680(.A(KEYINPUT118), .B(new_n675), .C1(new_n750), .C2(new_n652), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(new_n675), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n653), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n634), .A2(new_n643), .A3(new_n582), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n581), .B1(new_n646), .B2(new_n648), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n511), .B(new_n714), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n500), .A2(new_n501), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n438), .A2(new_n443), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n685), .A2(new_n877), .A3(new_n684), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n699), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n752), .A2(new_n769), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n755), .A2(new_n760), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n875), .A2(new_n704), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n680), .A2(new_n816), .A3(new_n697), .A4(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n707), .A2(new_n884), .B1(new_n772), .B2(new_n783), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n871), .A2(new_n881), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n866), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n729), .A2(new_n720), .A3(new_n721), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n746), .B1(new_n781), .B2(new_n782), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n692), .B(new_n705), .C1(new_n695), .C2(new_n696), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT120), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n718), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n733), .A2(new_n330), .A3(new_n684), .A4(new_n730), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n733), .B1(new_n707), .B2(new_n730), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n773), .A2(new_n708), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n888), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n732), .B2(new_n734), .ZN(new_n902));
  AOI22_X1  g716(.A1(new_n861), .A2(new_n772), .B1(new_n706), .B2(new_n707), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n901), .A2(KEYINPUT52), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT52), .B1(new_n901), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n887), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT53), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT52), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n895), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n773), .A2(new_n912), .A3(new_n708), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n773), .B2(new_n708), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n735), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n887), .B(new_n909), .C1(new_n906), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(KEYINPUT54), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n907), .A2(new_n909), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n887), .B(KEYINPUT53), .C1(new_n906), .C2(new_n916), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n865), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT124), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n865), .A2(new_n925), .A3(new_n918), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n503), .A2(new_n370), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n749), .A2(new_n746), .A3(new_n580), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n444), .A2(new_n668), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT49), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n744), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT117), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n718), .B(new_n725), .C1(new_n931), .C2(new_n744), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n937), .ZN(G75));
  XOR2_X1   g752(.A(KEYINPUT125), .B(KEYINPUT55), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n879), .B1(new_n748), .B2(new_n768), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(new_n752), .A3(new_n755), .A4(new_n760), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n749), .B(new_n651), .C1(new_n328), .C2(new_n329), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT118), .B1(new_n943), .B2(new_n675), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n653), .A2(new_n868), .A3(new_n869), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(new_n794), .A3(new_n796), .A4(new_n885), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n899), .A2(new_n900), .A3(new_n888), .ZN(new_n949));
  AOI21_X1  g763(.A(KEYINPUT121), .B1(new_n902), .B2(new_n903), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n910), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT52), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n920), .B1(new_n953), .B2(KEYINPUT53), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n655), .A3(new_n582), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n626), .A2(new_n628), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n632), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n645), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n955), .B2(new_n956), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n940), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n323), .B(new_n581), .C1(new_n919), .C2(new_n920), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n959), .B1(new_n964), .B2(KEYINPUT56), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n966), .A3(new_n939), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n370), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n963), .A2(new_n967), .A3(new_n969), .ZN(G51));
  XNOR2_X1  g784(.A(new_n954), .B(new_n921), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n575), .B(KEYINPUT57), .Z(new_n972));
  OAI22_X1  g786(.A1(new_n971), .A2(new_n972), .B1(new_n567), .B2(new_n564), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n954), .A2(new_n655), .A3(new_n811), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(G54));
  AND4_X1   g789(.A1(KEYINPUT58), .A2(new_n954), .A3(G475), .A4(new_n655), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n969), .B1(new_n976), .B2(new_n427), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n427), .B2(new_n976), .ZN(G60));
  NAND2_X1  g792(.A1(new_n658), .A2(new_n660), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT59), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n971), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n918), .A2(new_n922), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT60), .Z(new_n988));
  AND2_X1   g802(.A1(new_n954), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n375), .A2(new_n381), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n969), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n954), .A2(new_n691), .A3(new_n988), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n991), .B2(new_n993), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(G66));
  INV_X1    g810(.A(new_n947), .ZN(new_n997));
  NAND2_X1  g811(.A1(G224), .A2(G953), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n997), .A2(G953), .B1(new_n509), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(G898), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n957), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n999), .B(new_n1001), .ZN(G69));
  INV_X1    g816(.A(new_n831), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n735), .B1(new_n913), .B2(new_n914), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT126), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n914), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n903), .A2(new_n912), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n1006), .A2(new_n1007), .B1(new_n734), .B2(new_n732), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n1009), .A3(new_n831), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n815), .A2(new_n578), .A3(new_n710), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n393), .B(new_n889), .C1(new_n790), .C2(new_n791), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n794), .B(new_n796), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n839), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n370), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n370), .A2(G900), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(G953), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1022));
  OAI21_X1  g836(.A(KEYINPUT127), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n277), .A2(new_n285), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n422), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(G227), .A2(G900), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(G953), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1008), .A2(new_n726), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT62), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n750), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n669), .B1(new_n720), .B2(new_n875), .ZN(new_n1034));
  NOR4_X1   g848(.A1(new_n1033), .A2(new_n711), .A3(new_n776), .A4(new_n1034), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n839), .A2(new_n1003), .A3(new_n1035), .ZN(new_n1036));
  AND2_X1   g850(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  OR3_X1    g851(.A1(new_n1037), .A2(G953), .A3(new_n1026), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1027), .A2(new_n1029), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1024), .A2(G953), .A3(new_n1028), .A4(new_n1026), .ZN(new_n1040));
  AND2_X1   g854(.A1(new_n1039), .A2(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(new_n1037), .A2(new_n947), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT63), .Z(new_n1044));
  NAND2_X1  g858(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n321), .A2(new_n267), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n968), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1044), .B1(new_n1016), .B2(new_n997), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1048), .A2(new_n267), .A3(new_n321), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n289), .B1(new_n321), .B2(new_n266), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n908), .A2(new_n917), .A3(new_n1044), .A4(new_n1050), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(G57));
endmodule


