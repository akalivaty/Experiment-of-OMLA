//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT3), .A3(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n190), .B2(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(KEYINPUT80), .A3(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n192), .A2(new_n193), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n188), .A2(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n190), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT82), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G116), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT2), .B(G113), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT66), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT66), .B1(new_n204), .B2(new_n206), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT5), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n205), .A2(G119), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT5), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n209), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n197), .A2(new_n218), .A3(new_n200), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n202), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n203), .A2(G116), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n214), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n208), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n207), .A2(new_n208), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G101), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n234), .A3(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n220), .B1(new_n230), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G110), .B(G122), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n220), .B(new_n238), .C1(new_n230), .C2(new_n236), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n243), .A3(new_n239), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT64), .B1(new_n245), .B2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(G146), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n245), .B2(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n248), .A2(KEYINPUT65), .A3(G143), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .A4(new_n250), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n251), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n257), .A2(new_n258), .A3(new_n250), .A4(new_n264), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n255), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G224), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n270), .B(new_n272), .Z(new_n273));
  NAND3_X1  g087(.A1(new_n242), .A2(new_n244), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n238), .B(KEYINPUT8), .ZN(new_n275));
  INV_X1    g089(.A(new_n219), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n218), .B1(new_n197), .B2(new_n200), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n216), .B1(new_n215), .B2(new_n207), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n227), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n201), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n217), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n263), .A2(new_n269), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n272), .A2(new_n284), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n267), .A2(new_n268), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n262), .B(new_n286), .C1(new_n287), .C2(new_n255), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n241), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n274), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n274), .A2(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n274), .A2(new_n298), .A3(new_n292), .ZN(new_n299));
  INV_X1    g113(.A(new_n293), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT85), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n293), .B1(new_n296), .B2(KEYINPUT84), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT85), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n299), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n295), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT83), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n276), .A2(new_n277), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n254), .A2(new_n261), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n261), .A2(KEYINPUT81), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n257), .A2(new_n250), .A3(new_n258), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n253), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n197), .B(new_n200), .C1(KEYINPUT81), .C2(new_n261), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n309), .A2(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(G134), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n321), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n315), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n254), .A2(new_n330), .A3(new_n261), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n202), .A2(new_n219), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(KEYINPUT68), .A3(new_n325), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT68), .B1(new_n323), .B2(new_n325), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n233), .A2(new_n287), .A3(new_n235), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n313), .B2(new_n314), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n334), .A2(new_n339), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G140), .ZN(new_n344));
  INV_X1    g158(.A(G227), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT12), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n310), .B1(new_n202), .B2(new_n219), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n313), .A2(new_n314), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n338), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n328), .A2(new_n343), .A3(new_n348), .A4(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n342), .B(new_n340), .C1(new_n332), .C2(new_n333), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n354), .A2(new_n338), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n338), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(G469), .A2(G902), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n352), .B1(new_n354), .B2(new_n338), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n349), .B1(new_n315), .B2(new_n326), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n347), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n354), .A2(new_n338), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n343), .A2(new_n365), .A3(new_n348), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(G469), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(G221), .B1(new_n369), .B2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n306), .A2(new_n308), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT22), .B(G137), .ZN(new_n374));
  INV_X1    g188(.A(G953), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n375), .A2(G221), .A3(G234), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n374), .B(new_n376), .Z(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT75), .A2(G125), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G140), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT76), .B1(new_n381), .B2(G125), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(KEYINPUT75), .A3(G125), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT16), .A4(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n384), .A2(KEYINPUT77), .ZN(new_n389));
  OAI21_X1  g203(.A(G146), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G125), .B(G140), .Z(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G146), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT73), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n259), .A2(G119), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G110), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n203), .A2(G128), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n396), .B1(new_n203), .B2(G128), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n402), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT24), .B(G110), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n392), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n382), .A2(new_n383), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n386), .A3(KEYINPUT16), .A4(new_n380), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n384), .A2(new_n387), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n248), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n390), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n405), .A2(new_n406), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(G110), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n398), .B1(new_n395), .B2(new_n396), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n402), .ZN(new_n419));
  OAI21_X1  g233(.A(G110), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  AOI221_X4 g236(.A(KEYINPUT78), .B1(new_n390), .B2(new_n408), .C1(new_n413), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n422), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n390), .A2(new_n408), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n377), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n413), .A2(new_n422), .B1(new_n390), .B2(new_n408), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n377), .B1(new_n429), .B2(new_n424), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n428), .A2(new_n291), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n428), .A2(KEYINPUT25), .A3(new_n431), .A4(new_n291), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(G234), .B2(new_n291), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n373), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  AOI211_X1 g254(.A(KEYINPUT79), .B(new_n440), .C1(new_n434), .C2(new_n435), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n388), .A2(new_n389), .A3(G146), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n248), .B1(new_n410), .B2(new_n411), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n414), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n416), .B1(new_n415), .B2(G110), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n426), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n429), .A2(new_n424), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n430), .B1(new_n452), .B2(new_n377), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n438), .A2(G902), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n439), .A2(new_n441), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n457));
  INV_X1    g271(.A(new_n319), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n317), .A2(G137), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(new_n325), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n329), .A2(new_n461), .A3(new_n331), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n326), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n287), .A3(new_n335), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n230), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n287), .A2(new_n326), .B1(new_n461), .B2(new_n310), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n230), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n225), .A2(new_n227), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n326), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n267), .A2(new_n268), .ZN(new_n478));
  INV_X1    g292(.A(new_n312), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n479), .A2(new_n260), .B1(new_n251), .B2(new_n253), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n460), .A2(new_n325), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n477), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n476), .A2(new_n482), .A3(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n472), .A2(new_n466), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n469), .B1(KEYINPUT28), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(G237), .A2(G953), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT27), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT29), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT30), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n466), .ZN(new_n496));
  INV_X1    g310(.A(new_n490), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n457), .B1(new_n491), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(KEYINPUT28), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n490), .A3(new_n468), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n501), .A2(new_n457), .A3(new_n502), .A4(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(new_n462), .ZN(new_n504));
  INV_X1    g318(.A(new_n465), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n476), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n466), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n469), .B1(new_n507), .B2(KEYINPUT28), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n497), .A2(new_n502), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G472), .B1(new_n499), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT32), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT31), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n466), .A2(KEYINPUT70), .A3(new_n490), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n495), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT70), .B1(new_n466), .B2(new_n490), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n466), .A2(new_n490), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(KEYINPUT31), .A3(new_n495), .A4(new_n515), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n500), .A2(new_n468), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n497), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G472), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n518), .A2(new_n522), .B1(new_n524), .B2(new_n497), .ZN(new_n529));
  NOR4_X1   g343(.A1(new_n529), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n512), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n456), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(G143), .B1(new_n486), .B2(G214), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n486), .A2(G143), .A3(G214), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n390), .A2(new_n412), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n412), .A4(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(new_n535), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n542), .B2(new_n533), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n324), .A3(new_n535), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n541), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT18), .A2(G131), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n536), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n248), .B1(new_n409), .B2(new_n380), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n392), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(G113), .B(G122), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT86), .B(G104), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n549), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n549), .B2(new_n553), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n291), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT89), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n291), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(G475), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT13), .B1(new_n259), .B2(G143), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n317), .ZN(new_n566));
  XNOR2_X1  g380(.A(G128), .B(G143), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT90), .ZN(new_n569));
  INV_X1    g383(.A(G122), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(KEYINPUT90), .A2(G122), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n205), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n570), .A2(G116), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n190), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n573), .A2(G107), .A3(new_n574), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n568), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT14), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n574), .B(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G107), .B1(new_n580), .B2(new_n573), .ZN(new_n581));
  INV_X1    g395(.A(new_n577), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n567), .B(new_n317), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n369), .A2(new_n437), .A3(G953), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n578), .A2(new_n584), .ZN(new_n588));
  INV_X1    g402(.A(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n291), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n593), .B(new_n595), .Z(new_n596));
  NAND3_X1  g410(.A1(new_n549), .A2(new_n553), .A3(new_n557), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n543), .A2(new_n544), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n409), .A2(new_n380), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(KEYINPUT19), .B2(new_n391), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n598), .B1(new_n601), .B2(G146), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n553), .B1(new_n602), .B2(new_n443), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n556), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G475), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n291), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT20), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n597), .A2(new_n604), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT20), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n606), .A4(new_n291), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n564), .A2(new_n596), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G234), .ZN(new_n614));
  INV_X1    g428(.A(G237), .ZN(new_n615));
  OAI211_X1 g429(.A(G902), .B(G953), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT92), .Z(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT21), .B(G898), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n375), .A2(G952), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n614), .B2(new_n615), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n372), .A2(new_n532), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND2_X1  g440(.A1(new_n526), .A2(new_n527), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n529), .B2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT93), .A3(new_n628), .ZN(new_n629));
  OR3_X1    g443(.A1(new_n526), .A2(KEYINPUT93), .A3(new_n527), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n456), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n371), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n588), .B2(new_n589), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n592), .A2(new_n634), .B1(new_n586), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n594), .A2(G902), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(new_n594), .B2(new_n593), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n564), .B2(new_n612), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n293), .B1(new_n274), .B2(new_n292), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n308), .B1(new_n641), .B2(new_n294), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(new_n622), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n633), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND2_X1  g460(.A1(new_n564), .A2(new_n612), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n596), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  INV_X1    g463(.A(new_n308), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n622), .B(KEYINPUT94), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n650), .B(new_n651), .C1(new_n295), .C2(new_n640), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n596), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n564), .A3(new_n612), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT95), .B1(new_n656), .B2(new_n652), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n633), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT35), .B(G107), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  NOR2_X1   g475(.A1(new_n371), .A2(new_n308), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n304), .A2(new_n297), .A3(new_n299), .A4(new_n300), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n304), .B1(new_n303), .B2(new_n299), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n294), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n624), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT25), .B1(new_n453), .B2(new_n291), .ZN(new_n667));
  INV_X1    g481(.A(new_n435), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n438), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT79), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n436), .A2(new_n373), .A3(new_n438), .ZN(new_n671));
  INV_X1    g485(.A(new_n377), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n449), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n454), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n670), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n631), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n666), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(new_n371), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n531), .A2(new_n676), .A3(new_n681), .A4(new_n642), .ZN(new_n682));
  INV_X1    g496(.A(new_n621), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n683), .B1(new_n617), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n656), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XNOR2_X1  g502(.A(new_n665), .B(KEYINPUT38), .ZN(new_n689));
  INV_X1    g503(.A(new_n647), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n676), .A2(new_n690), .A3(new_n596), .A4(new_n308), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n521), .A2(new_n495), .A3(new_n515), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n507), .A2(new_n497), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n528), .B2(new_n530), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT96), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n699), .B(new_n696), .C1(new_n528), .C2(new_n530), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT97), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n689), .A2(new_n701), .A3(KEYINPUT97), .A4(new_n691), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n685), .B(new_n704), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n681), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT40), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT99), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n689), .A2(new_n691), .ZN(new_n711));
  INV_X1    g525(.A(new_n701), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n714), .A3(new_n703), .A4(new_n707), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n245), .ZN(G45));
  AOI211_X1 g531(.A(new_n685), .B(new_n638), .C1(new_n564), .C2(new_n612), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n682), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(new_n456), .A2(new_n531), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n362), .A2(new_n363), .A3(new_n347), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n348), .B1(new_n343), .B2(new_n365), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n291), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n360), .A3(new_n370), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n643), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n658), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  NOR3_X1   g546(.A1(new_n613), .A2(new_n726), .A3(new_n623), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n531), .A3(new_n642), .A4(new_n676), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  AND3_X1   g549(.A1(new_n647), .A2(new_n655), .A3(new_n642), .ZN(new_n736));
  INV_X1    g550(.A(new_n726), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n651), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n508), .A2(new_n490), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n523), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n527), .A2(new_n291), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n628), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n456), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n570), .ZN(G24));
  NOR2_X1   g560(.A1(new_n439), .A2(new_n441), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n742), .B1(new_n747), .B2(new_n675), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT100), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n650), .B1(new_n295), .B2(new_n640), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n726), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n749), .A3(new_n718), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n676), .A2(new_n718), .A3(new_n743), .A4(new_n751), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT100), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  OAI211_X1 g570(.A(new_n294), .B(new_n650), .C1(new_n663), .C2(new_n664), .ZN(new_n757));
  INV_X1    g571(.A(new_n370), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n364), .A2(new_n366), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT102), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n364), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(G469), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n361), .B(KEYINPUT101), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n358), .B2(new_n359), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n758), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT103), .B1(new_n757), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT103), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n306), .A2(new_n770), .A3(new_n650), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n718), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT42), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(KEYINPUT104), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n774), .A2(KEYINPUT104), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n532), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n721), .B1(new_n769), .B2(new_n771), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n778), .B2(new_n775), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n686), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  INV_X1    g597(.A(new_n638), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n690), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT43), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n676), .A2(new_n630), .A3(new_n629), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n757), .B1(new_n788), .B2(KEYINPUT44), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n760), .A2(KEYINPUT45), .A3(new_n762), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n359), .B1(new_n759), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n765), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT105), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n793), .A2(new_n794), .A3(KEYINPUT46), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n724), .A2(G469), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n793), .B2(KEYINPUT46), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n370), .A3(new_n705), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n789), .B(new_n800), .C1(KEYINPUT44), .C2(new_n788), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(new_n757), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n718), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n804), .A2(new_n531), .A3(new_n456), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n370), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(KEYINPUT106), .A3(new_n370), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT107), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(KEYINPUT107), .A3(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(KEYINPUT107), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n809), .A4(new_n811), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n805), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT108), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND2_X1  g633(.A1(new_n712), .A2(new_n456), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n725), .A2(new_n360), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n308), .B(new_n758), .C1(new_n821), .C2(KEYINPUT49), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(KEYINPUT49), .B2(new_n821), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n820), .A2(new_n689), .A3(new_n785), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT109), .Z(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n727), .B1(new_n643), .B2(new_n658), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT110), .B1(new_n648), .B2(new_n639), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n656), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n631), .A2(new_n456), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n372), .A3(new_n832), .A4(new_n651), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n833), .A3(new_n734), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n738), .A2(new_n744), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n678), .A2(new_n835), .A3(new_n625), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n752), .A2(new_n754), .B1(new_n682), .B2(new_n686), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n767), .A2(new_n655), .A3(new_n647), .A4(new_n642), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n698), .B2(new_n700), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT112), .B1(new_n676), .B2(new_n685), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  INV_X1    g656(.A(new_n685), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n747), .A2(new_n842), .A3(new_n675), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n840), .A2(new_n845), .B1(new_n682), .B2(new_n718), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n838), .A2(new_n846), .A3(KEYINPUT52), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(new_n838), .B2(new_n846), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n780), .B(new_n837), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n748), .A2(new_n718), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n531), .A2(new_n676), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n367), .A2(new_n361), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n370), .B(new_n843), .C1(new_n797), .C2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n757), .A2(new_n613), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n772), .A2(new_n850), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n856), .A2(new_n782), .A3(KEYINPUT111), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT111), .B1(new_n856), .B2(new_n782), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n826), .B1(new_n849), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n666), .B1(new_n721), .B2(new_n677), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n745), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n734), .A3(new_n827), .A4(new_n833), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n779), .A3(new_n777), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n782), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n856), .A2(new_n782), .A3(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n838), .A2(new_n846), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n838), .A2(new_n846), .A3(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n864), .A2(new_n869), .A3(new_n874), .A4(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n860), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n860), .A2(new_n875), .A3(KEYINPUT54), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n786), .A2(new_n621), .A3(new_n744), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n689), .A2(new_n650), .A3(new_n726), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT50), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n803), .A2(new_n683), .A3(new_n737), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n786), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n748), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT114), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n820), .A2(new_n647), .A3(new_n784), .A4(new_n886), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n885), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n813), .A2(new_n815), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n821), .A2(new_n370), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n803), .B(new_n882), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n881), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n882), .A2(new_n751), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n620), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n887), .A2(new_n532), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT48), .Z(new_n901));
  NOR2_X1   g715(.A1(new_n820), .A2(new_n886), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n899), .B(new_n901), .C1(new_n639), .C2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n895), .B2(new_n896), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n880), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n825), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n375), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n291), .B1(new_n860), .B2(new_n875), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT56), .B1(new_n910), .B2(G210), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n242), .A2(new_n244), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n273), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n909), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(KEYINPUT116), .A3(G210), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT116), .B1(new_n910), .B2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n917), .B2(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n764), .B(KEYINPUT57), .Z(new_n923));
  NAND3_X1  g737(.A1(new_n878), .A2(new_n879), .A3(new_n923), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n924), .A2(KEYINPUT117), .B1(new_n357), .B2(new_n353), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(KEYINPUT117), .B2(new_n924), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n910), .A2(new_n790), .A3(new_n792), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n908), .B1(new_n926), .B2(new_n927), .ZN(G54));
  AND2_X1   g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n910), .A2(new_n609), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n609), .B1(new_n910), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n908), .ZN(G60));
  XNOR2_X1  g746(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n594), .A2(new_n291), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n880), .A2(new_n636), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n636), .B1(new_n880), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n908), .ZN(G63));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  XNOR2_X1  g753(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n437), .A2(new_n291), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n860), .B2(new_n875), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n944), .A2(KEYINPUT120), .A3(new_n674), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT120), .B1(new_n944), .B2(new_n674), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT121), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n909), .B1(new_n944), .B2(new_n453), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT122), .B(new_n909), .C1(new_n944), .C2(new_n453), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n939), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n954));
  OAI221_X1 g768(.A(new_n954), .B1(KEYINPUT121), .B2(KEYINPUT61), .C1(new_n946), .C2(new_n945), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n618), .B2(new_n271), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n837), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n912), .B1(G898), .B2(new_n375), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  AND2_X1   g774(.A1(new_n838), .A2(new_n719), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n709), .A2(new_n715), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT62), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n706), .A2(new_n757), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n831), .A2(new_n964), .A3(new_n532), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n801), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n805), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n817), .B1(new_n892), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g782(.A(KEYINPUT108), .B(new_n805), .C1(new_n813), .C2(new_n815), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n375), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n492), .A2(new_n494), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT123), .Z(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(new_n601), .Z(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT124), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n345), .B2(new_n684), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT125), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n800), .A2(new_n532), .A3(new_n736), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n782), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n780), .A2(new_n801), .A3(new_n980), .A4(new_n961), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n968), .B2(new_n969), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n375), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n684), .A2(G953), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n974), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n976), .B(new_n978), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n978), .ZN(new_n988));
  INV_X1    g802(.A(new_n975), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n962), .B(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n818), .A3(new_n966), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n989), .B1(new_n992), .B2(new_n375), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n986), .B1(new_n983), .B2(new_n984), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n987), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(new_n496), .A2(new_n490), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n991), .A2(new_n818), .A3(new_n837), .A4(new_n966), .ZN(new_n998));
  XNOR2_X1  g812(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n527), .A2(new_n291), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n999), .B(new_n1000), .Z(new_n1001));
  AOI21_X1  g815(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g818(.A(KEYINPUT127), .B(new_n997), .C1(new_n998), .C2(new_n1001), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1001), .B1(new_n982), .B2(new_n863), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1006), .A2(new_n497), .A3(new_n466), .A4(new_n495), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1001), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n693), .B2(new_n498), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n908), .B1(new_n876), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n1004), .A2(new_n1005), .A3(new_n1011), .ZN(G57));
endmodule


