//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n198), .A2(new_n190), .A3(new_n192), .A4(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n197), .A3(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n198), .A2(new_n189), .A3(G146), .A4(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G134), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n209), .A3(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT30), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n218), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n195), .A2(KEYINPUT0), .A3(new_n196), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n194), .A2(new_n197), .A3(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n217), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n215), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n230), .A3(new_n214), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n203), .A3(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n190), .A2(new_n192), .A3(new_n196), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n196), .B1(new_n190), .B2(new_n192), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n223), .B1(new_n235), .B2(KEYINPUT0), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT67), .B1(new_n236), .B2(new_n222), .ZN(new_n237));
  AND4_X1   g051(.A1(KEYINPUT67), .A2(new_n222), .A3(new_n224), .A4(new_n225), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n228), .B1(new_n239), .B2(KEYINPUT30), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT2), .B(G113), .Z(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n241), .A2(KEYINPUT66), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT66), .B1(new_n241), .B2(new_n242), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(new_n241), .B2(new_n242), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n188), .B1(new_n240), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G237), .ZN(new_n248));
  INV_X1    g062(.A(G953), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G210), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n226), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n222), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n212), .A2(new_n230), .A3(new_n214), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n230), .B1(new_n212), .B2(new_n214), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n256), .A2(new_n257), .B1(new_n260), .B2(new_n203), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n246), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(new_n257), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n217), .B1(new_n263), .B2(new_n232), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT69), .B(new_n245), .C1(new_n264), .C2(new_n228), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n247), .A2(new_n254), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n232), .A2(new_n246), .A3(new_n226), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT28), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT71), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n216), .A2(new_n226), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n245), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n245), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n262), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n254), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n267), .A2(new_n268), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n187), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n240), .A2(new_n188), .A3(new_n246), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n227), .B1(new_n261), .B2(new_n217), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT69), .B1(new_n287), .B2(new_n245), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n254), .A4(new_n262), .ZN(new_n291));
  INV_X1    g105(.A(new_n254), .ZN(new_n292));
  INV_X1    g106(.A(new_n280), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n272), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n283), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(KEYINPUT72), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n283), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(new_n187), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n239), .B(new_n246), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(new_n270), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT29), .B1(new_n303), .B2(new_n272), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n273), .A2(new_n280), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n304), .B(new_n254), .C1(KEYINPUT29), .C2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n289), .A2(new_n292), .A3(new_n262), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n306), .B(new_n307), .C1(KEYINPUT29), .C2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n298), .A2(new_n301), .B1(G472), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(KEYINPUT73), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n196), .A2(G119), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n319), .B2(G110), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n314), .A2(G128), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT24), .B(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT76), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n315), .A2(new_n326), .A3(new_n327), .A4(new_n318), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT16), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n330), .A3(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT74), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n334), .B2(new_n337), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(new_n340), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n334), .A2(G146), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT78), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n329), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n319), .A2(G110), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n336), .B2(new_n340), .ZN(new_n348));
  INV_X1    g162(.A(new_n341), .ZN(new_n349));
  OAI221_X1 g163(.A(new_n347), .B1(new_n322), .B2(new_n323), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n350), .A3(KEYINPUT80), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(G137), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n354), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n352), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n363), .C2(G902), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(G234), .B2(new_n307), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n362), .A2(new_n307), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n366), .A2(G902), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n362), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n310), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(KEYINPUT3), .A2(G107), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT83), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G104), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT3), .A2(G107), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n380), .A2(new_n382), .ZN(new_n392));
  INV_X1    g206(.A(new_n378), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n386), .A2(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(new_n251), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT84), .B(G101), .C1(new_n383), .C2(new_n388), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n391), .A2(new_n396), .A3(KEYINPUT4), .A4(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(G101), .C1(new_n383), .C2(new_n388), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT83), .B(G104), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n386), .B(new_n387), .C1(new_n403), .C2(new_n378), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(KEYINPUT85), .A3(new_n399), .A4(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n245), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n314), .A2(G116), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n408), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT88), .B1(new_n408), .B2(KEYINPUT5), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n409), .A2(new_n410), .A3(G113), .A4(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n243), .B2(new_n244), .ZN(new_n413));
  NAND2_X1  g227(.A1(G104), .A2(G107), .ZN(new_n414));
  OAI211_X1 g228(.A(G101), .B(new_n414), .C1(new_n403), .C2(G107), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n396), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G122), .Z(new_n420));
  AND4_X1   g234(.A1(KEYINPUT90), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n407), .B2(new_n417), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT90), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n419), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n413), .A2(new_n416), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n383), .A2(new_n388), .A3(G101), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n390), .B2(new_n389), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n430), .A2(new_n431), .B1(new_n402), .B2(new_n405), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n428), .B1(new_n432), .B2(new_n245), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT89), .B1(new_n433), .B2(new_n422), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n422), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n236), .A2(G125), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n203), .A2(new_n332), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G224), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(G953), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n439), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n425), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n420), .B(KEYINPUT8), .Z(new_n444));
  AND2_X1   g258(.A1(new_n413), .A2(new_n416), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n428), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(new_n440), .B2(G953), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n447), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n435), .A2(new_n446), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n450), .A2(new_n307), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n443), .A2(new_n453), .A3(new_n451), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G116), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G122), .ZN(new_n465));
  INV_X1    g279(.A(G122), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G116), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n468), .B(KEYINPUT97), .Z(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n385), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n196), .A2(G143), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n189), .A2(G128), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(new_n205), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n465), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT99), .B1(new_n465), .B2(KEYINPUT14), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(KEYINPUT14), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n475), .A2(new_n467), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G107), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT100), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT100), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n470), .A2(new_n482), .A3(new_n474), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(new_n205), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n471), .A2(KEYINPUT13), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT98), .ZN(new_n487));
  INV_X1    g301(.A(new_n472), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n471), .B2(KEYINPUT13), .ZN(new_n489));
  OAI21_X1  g303(.A(G134), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n470), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n469), .A2(new_n385), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n485), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(KEYINPUT9), .B(G234), .Z(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(new_n365), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n484), .A2(new_n493), .A3(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n463), .B1(new_n501), .B2(new_n307), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n484), .A2(new_n493), .A3(new_n497), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n497), .B1(new_n484), .B2(new_n493), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n307), .B(new_n463), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n248), .A2(new_n249), .A3(G214), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(G143), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT92), .B(G143), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G131), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(KEYINPUT93), .A3(G131), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT17), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n513), .A2(G131), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n516), .A2(new_n520), .A3(new_n521), .A4(new_n517), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT94), .B1(new_n349), .B2(new_n348), .ZN(new_n523));
  INV_X1    g337(.A(new_n348), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n341), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n519), .A2(new_n522), .A3(new_n523), .A4(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n379), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n345), .B1(new_n191), .B2(new_n335), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n513), .A2(KEYINPUT18), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n513), .A2(KEYINPUT18), .A3(G131), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n530), .A2(new_n520), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n529), .B1(new_n527), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n307), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT96), .B(G475), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n516), .A2(new_n520), .A3(new_n517), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n334), .B(KEYINPUT19), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n343), .B(new_n540), .C1(G146), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  INV_X1    g357(.A(new_n529), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n527), .A2(new_n529), .A3(new_n533), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT95), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n539), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  AOI211_X1 g365(.A(KEYINPUT20), .B(new_n549), .C1(new_n545), .C2(new_n546), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n538), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G952), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G953), .ZN(new_n555));
  NAND2_X1  g369(.A1(G234), .A2(G237), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT21), .B(G898), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(G902), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n508), .A2(new_n553), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n460), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n458), .B1(new_n457), .B2(new_n459), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n249), .A2(G227), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT82), .ZN(new_n569));
  XNOR2_X1  g383(.A(G110), .B(G140), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n432), .A2(new_n236), .ZN(new_n572));
  INV_X1    g386(.A(new_n416), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT1), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n201), .B1(new_n574), .B2(new_n190), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n203), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n572), .A2(new_n582), .A3(new_n578), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n222), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n222), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n572), .A2(new_n585), .A3(new_n578), .A4(new_n579), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n571), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n571), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n416), .A2(new_n202), .A3(new_n201), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(KEYINPUT86), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n585), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n576), .A2(KEYINPUT86), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT12), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n594), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n588), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n567), .B(new_n307), .C1(new_n587), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G469), .A2(G902), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n584), .A2(new_n586), .A3(new_n571), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n580), .A2(new_n222), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n571), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n599), .B(new_n600), .C1(new_n604), .C2(new_n567), .ZN(new_n605));
  OAI21_X1  g419(.A(G221), .B1(new_n496), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n565), .A2(new_n566), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n377), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  NOR2_X1   g424(.A1(new_n376), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n296), .A2(new_n307), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT101), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n615), .A3(G472), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n611), .A2(new_n299), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT102), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n614), .A2(new_n616), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n299), .A4(new_n611), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n456), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n443), .A2(new_n451), .A3(KEYINPUT103), .A4(new_n453), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n452), .B2(new_n454), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT104), .B(new_n453), .C1(new_n443), .C2(new_n451), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n623), .B(new_n624), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n459), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n618), .A2(new_n621), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n503), .A2(new_n504), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT33), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n501), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n633), .A2(new_n635), .A3(G478), .A4(new_n307), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT105), .B(G478), .Z(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n632), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n553), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n563), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n631), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n553), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n563), .B(KEYINPUT106), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n645), .A2(new_n508), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n631), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n351), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n374), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n373), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n608), .A2(new_n619), .A3(new_n299), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n558), .B1(new_n562), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n553), .A2(new_n507), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n626), .A2(new_n627), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n623), .A2(new_n624), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n459), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n628), .A2(KEYINPUT108), .A3(new_n459), .A4(new_n661), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n309), .A2(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT32), .B1(new_n296), .B2(new_n283), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n301), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n607), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n668), .A2(new_n674), .A3(new_n675), .A4(new_n654), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT109), .ZN(new_n677));
  INV_X1    g491(.A(new_n654), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n298), .A2(new_n301), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n669), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n675), .A4(new_n668), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  NAND2_X1  g498(.A1(new_n289), .A2(new_n262), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n254), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n302), .B2(new_n292), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n298), .A2(new_n301), .B1(G472), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n660), .B(KEYINPUT39), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n607), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n457), .B(KEYINPUT38), .Z(new_n694));
  NOR3_X1   g508(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n508), .A2(new_n553), .A3(new_n459), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n654), .B(new_n698), .C1(new_n692), .C2(new_n691), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n189), .ZN(G45));
  NOR2_X1   g514(.A1(new_n640), .A2(new_n660), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n459), .A3(new_n628), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n310), .A2(new_n607), .A3(new_n678), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n191), .ZN(G48));
  INV_X1    g518(.A(new_n376), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n307), .B1(new_n587), .B2(new_n598), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G469), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n707), .A2(new_n606), .A3(new_n599), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n629), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n674), .A2(new_n705), .A3(new_n641), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND4_X1  g527(.A1(new_n674), .A2(new_n647), .A3(new_n705), .A4(new_n710), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NAND4_X1  g529(.A1(new_n674), .A2(new_n564), .A3(new_n654), .A4(new_n710), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  INV_X1    g531(.A(new_n613), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n267), .A2(new_n268), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n292), .B1(new_n303), .B2(new_n272), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n284), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n718), .A2(new_n376), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n697), .A2(new_n628), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n646), .A3(new_n708), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(G122), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G24));
  NOR3_X1   g540(.A1(new_n678), .A2(new_n718), .A3(new_n721), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n701), .A3(new_n710), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n332), .ZN(G27));
  NAND3_X1  g543(.A1(new_n669), .A2(new_n285), .A3(new_n297), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n705), .ZN(new_n731));
  INV_X1    g545(.A(new_n459), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n457), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n675), .A2(new_n701), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT42), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n674), .A2(new_n705), .A3(new_n675), .A4(new_n733), .ZN(new_n736));
  OR3_X1    g550(.A1(new_n640), .A2(KEYINPUT42), .A3(new_n660), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n211), .ZN(G33));
  INV_X1    g553(.A(new_n661), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n205), .ZN(G36));
  INV_X1    g556(.A(new_n639), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n553), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(KEYINPUT43), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(KEYINPUT43), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n744), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n747), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n678), .B1(new_n619), .B2(new_n299), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT44), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(new_n733), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(KEYINPUT112), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n751), .A2(new_n752), .ZN(new_n758));
  AOI211_X1 g572(.A(new_n755), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n604), .B(KEYINPUT45), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n760), .B2(G902), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n599), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n606), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n690), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G137), .ZN(G39));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n765), .B1(new_n769), .B2(KEYINPUT47), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n772));
  MUX2_X1   g586(.A(new_n770), .B(new_n765), .S(new_n772), .Z(new_n773));
  NAND4_X1  g587(.A1(new_n310), .A2(new_n376), .A3(new_n701), .A4(new_n733), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT114), .Z(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n330), .ZN(G42));
  NAND2_X1  g591(.A1(new_n554), .A2(new_n249), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n508), .A2(new_n553), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n680), .A2(new_n675), .A3(new_n779), .A4(new_n733), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n780), .B2(new_n660), .ZN(new_n781));
  INV_X1    g595(.A(new_n733), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n310), .A2(new_n607), .A3(new_n678), .A4(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  INV_X1    g598(.A(new_n660), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n779), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n640), .B1(new_n507), .B2(new_n553), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n460), .A3(new_n646), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n566), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n618), .A2(new_n621), .A3(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n791), .A2(new_n609), .A3(new_n655), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n734), .A2(new_n718), .A3(new_n678), .A4(new_n721), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n741), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n787), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n711), .A2(new_n714), .A3(new_n716), .A4(new_n724), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n738), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n703), .ZN(new_n800));
  INV_X1    g614(.A(new_n728), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n689), .A2(new_n607), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n678), .A3(new_n785), .A4(new_n723), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n683), .A2(new_n800), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n728), .B1(new_n677), .B2(new_n682), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(KEYINPUT52), .A3(new_n800), .A4(new_n803), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n804), .B2(new_n805), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n799), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n787), .A2(new_n797), .A3(new_n792), .A4(new_n794), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n728), .B(new_n703), .C1(new_n677), .C2(new_n682), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(new_n814), .B2(new_n803), .ZN(new_n815));
  AND4_X1   g629(.A1(KEYINPUT52), .A2(new_n807), .A3(new_n800), .A4(new_n803), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n812), .A2(new_n818), .A3(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n812), .A2(new_n818), .A3(new_n821), .A4(KEYINPUT54), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n787), .A2(new_n792), .A3(new_n794), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n798), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n795), .A2(KEYINPUT118), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n826), .B(new_n827), .C1(new_n811), .C2(new_n809), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n828), .B2(KEYINPUT53), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n820), .B(new_n822), .C1(KEYINPUT54), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n557), .B1(new_n748), .B2(new_n750), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n709), .A2(new_n782), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n731), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT48), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n705), .A2(new_n689), .A3(new_n558), .A4(new_n832), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n553), .A3(new_n639), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n722), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n554), .B(G953), .C1(new_n840), .C2(new_n710), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT121), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n707), .A2(new_n599), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n773), .B1(new_n606), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n733), .A3(new_n840), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n694), .A2(new_n732), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n831), .A2(new_n708), .A3(new_n722), .A4(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n727), .A2(new_n833), .B1(new_n848), .B2(KEYINPUT50), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n837), .A2(new_n645), .A3(new_n743), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n849), .B(new_n850), .C1(KEYINPUT50), .C2(new_n848), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT51), .B(new_n846), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n773), .A2(KEYINPUT119), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n844), .A2(new_n606), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n773), .B2(KEYINPUT119), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n782), .B(new_n839), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n851), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n843), .B(new_n855), .C1(new_n860), .C2(KEYINPUT51), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n778), .B1(new_n830), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n749), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n844), .A2(KEYINPUT49), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n705), .A2(new_n864), .A3(new_n694), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n459), .A3(new_n606), .A4(new_n689), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT122), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n862), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(G75));
  NAND2_X1  g686(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n873));
  INV_X1    g687(.A(new_n823), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n307), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G210), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n425), .A2(new_n436), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n442), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n877), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n877), .B2(new_n878), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n249), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(new_n600), .A2(KEYINPUT57), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n600), .A2(KEYINPUT57), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n587), .B2(new_n598), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n876), .A2(G469), .A3(new_n760), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n884), .B1(new_n891), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n546), .A3(new_n545), .ZN(new_n895));
  INV_X1    g709(.A(new_n884), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .A4(new_n547), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G60));
  AND2_X1   g712(.A1(new_n633), .A2(new_n635), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT59), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n899), .B(new_n901), .C1(new_n888), .C2(new_n889), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n830), .B2(new_n901), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n884), .A3(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT124), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n875), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n884), .B1(new_n910), .B2(new_n363), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n875), .A2(new_n909), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n652), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(new_n913), .C1(KEYINPUT125), .C2(KEYINPUT61), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n913), .B(new_n896), .C1(new_n362), .C2(new_n912), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT61), .B1(new_n913), .B2(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n560), .B2(new_n440), .ZN(new_n919));
  INV_X1    g733(.A(new_n792), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n796), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n921), .B2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n879), .B1(G898), .B2(new_n249), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G69));
  XOR2_X1   g738(.A(new_n541), .B(KEYINPUT126), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n240), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n249), .B1(G227), .B2(G900), .ZN(new_n927));
  INV_X1    g741(.A(new_n814), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n928), .A2(new_n699), .ZN(new_n929));
  XOR2_X1   g743(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n930));
  OR2_X1    g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n776), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n377), .A2(new_n691), .A3(new_n733), .A4(new_n788), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n933), .A2(new_n767), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI211_X1 g750(.A(new_n926), .B(new_n927), .C1(new_n936), .C2(new_n249), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n834), .A2(new_n723), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n759), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n738), .B1(new_n939), .B2(new_n766), .ZN(new_n940));
  INV_X1    g754(.A(new_n741), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n776), .A2(new_n928), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n940), .A2(new_n249), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n659), .B2(G227), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n937), .B1(new_n945), .B2(new_n926), .ZN(G72));
  NAND2_X1  g760(.A1(new_n686), .A2(new_n308), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  OAI21_X1  g764(.A(new_n896), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n818), .A2(new_n812), .A3(new_n950), .A4(new_n948), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n953), .A2(new_n308), .B1(new_n936), .B2(new_n686), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n951), .B(new_n952), .C1(new_n954), .C2(new_n921), .ZN(G57));
endmodule


