//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT81), .Z(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT74), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT2), .B1(new_n206), .B2(new_n208), .ZN(new_n217));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n214), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n211), .A2(new_n216), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G211gat), .A2(G218gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT22), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n223), .A3(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n222), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n210), .B(new_n212), .C1(new_n215), .C2(new_n213), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n215), .A2(new_n218), .ZN(new_n238));
  XNOR2_X1  g037(.A(G141gat), .B(G148gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT2), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n240), .A3(new_n235), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n232), .B1(new_n241), .B2(new_n233), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n204), .B1(new_n236), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(new_n234), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(KEYINPUT82), .A3(new_n233), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n222), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n242), .A2(new_n203), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n202), .B(new_n243), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(KEYINPUT83), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(KEYINPUT83), .ZN(new_n251));
  XNOR2_X1  g050(.A(G78gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT31), .B(G50gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  OAI21_X1  g053(.A(new_n243), .B1(new_n247), .B2(new_n248), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(G22gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n250), .A2(new_n256), .A3(KEYINPUT84), .A4(new_n251), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(G22gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n249), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n254), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT23), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n268), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT64), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G183gat), .A2(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT25), .ZN(new_n278));
  INV_X1    g077(.A(G169gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n270), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n272), .A2(new_n277), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n274), .A2(new_n273), .B1(new_n287), .B2(G190gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n268), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n289), .A3(new_n270), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n278), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT27), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n294), .B(KEYINPUT28), .C1(new_n299), .C2(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n281), .A2(KEYINPUT26), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT26), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n279), .A3(new_n280), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n270), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT27), .B(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n294), .A2(KEYINPUT28), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n307), .B2(KEYINPUT65), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n300), .A2(new_n274), .A3(new_n304), .A4(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n292), .A2(new_n293), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n293), .B1(new_n292), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n267), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n309), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n306), .B1(new_n305), .B2(new_n308), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n304), .A2(new_n274), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n316), .A2(new_n317), .B1(new_n286), .B2(new_n291), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT71), .B(new_n266), .C1(new_n318), .C2(KEYINPUT29), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n292), .B2(new_n310), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(new_n267), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n232), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT73), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n311), .A2(new_n312), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n266), .A2(new_n233), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n292), .A2(new_n310), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n329), .A2(new_n330), .B1(new_n266), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n232), .ZN(new_n333));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  NAND4_X1  g135(.A1(new_n326), .A2(new_n328), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(new_n328), .A3(new_n333), .ZN(new_n340));
  INV_X1    g139(.A(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n325), .A2(KEYINPUT73), .B1(new_n332), .B2(new_n232), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(KEYINPUT30), .A3(new_n328), .A4(new_n336), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G225gat), .A2(G233gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n346), .B(KEYINPUT75), .Z(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G113gat), .ZN(new_n349));
  INV_X1    g148(.A(G113gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G120gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n351), .A3(KEYINPUT66), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n348), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  XNOR2_X1  g153(.A(G127gat), .B(G134gat), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G127gat), .B(G134gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G113gat), .B(G120gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(KEYINPUT1), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n221), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n237), .A2(new_n240), .B1(new_n356), .B2(new_n359), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n347), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n360), .A3(new_n241), .ZN(new_n366));
  INV_X1    g165(.A(new_n360), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n360), .B2(new_n221), .ZN(new_n370));
  INV_X1    g169(.A(new_n347), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(new_n368), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n373), .B(new_n347), .C1(new_n361), .C2(new_n362), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n364), .A2(new_n372), .A3(KEYINPUT5), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n370), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n360), .A2(new_n221), .A3(new_n369), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT79), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(new_n370), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n347), .A2(KEYINPUT5), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n378), .A2(new_n380), .A3(new_n366), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(new_n380), .A3(new_n366), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n347), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n361), .A2(new_n362), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n393), .B(KEYINPUT39), .C1(new_n347), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n396), .A3(new_n347), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n397), .A2(KEYINPUT85), .A3(new_n389), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT85), .B1(new_n397), .B2(new_n389), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n395), .B(KEYINPUT40), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT40), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n345), .A2(new_n391), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n326), .A2(new_n405), .A3(new_n328), .A4(new_n333), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT86), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n343), .A2(new_n408), .A3(new_n405), .A4(new_n328), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n405), .B1(new_n332), .B2(new_n324), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n323), .A2(new_n232), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT38), .B(new_n336), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n375), .A2(new_n382), .A3(new_n389), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n389), .B1(new_n375), .B2(new_n382), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n418), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT87), .B1(new_n418), .B2(KEYINPUT6), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n337), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT38), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n336), .B1(new_n340), .B2(KEYINPUT37), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n410), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n265), .B(new_n404), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(KEYINPUT6), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n339), .A2(new_n430), .A3(new_n342), .A4(new_n344), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n338), .A2(new_n337), .B1(new_n417), .B2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n342), .A4(new_n344), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n259), .A2(new_n260), .B1(new_n263), .B2(new_n254), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  XOR2_X1   g238(.A(G15gat), .B(G43gat), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT69), .ZN(new_n441));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n331), .A2(new_n367), .ZN(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n292), .A2(new_n360), .A3(new_n310), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT67), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n444), .A2(new_n450), .A3(new_n446), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n443), .B1(new_n452), .B2(KEYINPUT32), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT68), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n456));
  AOI211_X1 g255(.A(new_n456), .B(KEYINPUT33), .C1(new_n449), .C2(new_n451), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n444), .A2(new_n447), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n445), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT34), .B1(new_n446), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n460), .B(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n452), .B(KEYINPUT32), .C1(new_n454), .C2(new_n443), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n458), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n439), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(new_n463), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT36), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n428), .A2(new_n438), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n465), .A2(new_n466), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n432), .A2(new_n435), .A3(new_n475), .A4(new_n265), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n437), .A2(new_n465), .A3(new_n466), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT35), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n421), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n345), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n476), .A2(KEYINPUT35), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(G197gat), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT11), .B(G169gat), .Z(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n486), .B(KEYINPUT12), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G29gat), .ZN(new_n489));
  INV_X1    g288(.A(G36gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT14), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n494), .A2(KEYINPUT88), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G43gat), .B(G50gat), .Z(new_n498));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n494), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n498), .A2(new_n499), .B1(G29gat), .B2(G36gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n501), .A2(new_n502), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(KEYINPUT17), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(G1gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT16), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(G1gat), .B2(new_n512), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(G8gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(G8gat), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n507), .B2(new_n509), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n511), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n508), .A2(new_n510), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n522), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n527), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n510), .A3(new_n508), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n529), .B(KEYINPUT13), .Z(new_n535));
  AOI22_X1  g334(.A1(new_n530), .A2(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n522), .A2(new_n528), .A3(KEYINPUT18), .A4(new_n529), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n488), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n488), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n482), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(G57gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G64gat), .ZN(new_n545));
  INV_X1    g344(.A(G64gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G57gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n545), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT93), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(G71gat), .A2(G78gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n555), .B2(new_n554), .ZN(new_n557));
  INV_X1    g356(.A(new_n547), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n546), .A2(G57gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT9), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT21), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G127gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n532), .B1(new_n563), .B2(new_n562), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  INV_X1    g375(.A(G92gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT7), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n575), .B(new_n581), .C1(new_n576), .C2(new_n577), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n583), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n580), .A2(new_n588), .A3(new_n582), .A4(new_n584), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT95), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n523), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n511), .A2(new_n521), .A3(new_n591), .ZN(new_n595));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n594), .B2(new_n595), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n562), .A2(new_n590), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n553), .A2(new_n587), .A3(new_n561), .A4(new_n589), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n591), .A2(new_n613), .A3(new_n562), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT96), .B1(new_n609), .B2(KEYINPUT10), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT96), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n616), .A3(new_n613), .A4(new_n608), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n610), .B(KEYINPUT97), .Z(new_n619));
  OAI21_X1  g418(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n612), .B(new_n623), .C1(new_n618), .C2(new_n611), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g426(.A1(new_n574), .A2(new_n606), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n543), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n430), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n513), .ZN(G1324gat));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n345), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT16), .B(G8gat), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT42), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n635), .A2(new_n636), .B1(G8gat), .B2(new_n633), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(G1325gat));
  AND3_X1   g437(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT98), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT98), .B1(new_n467), .B2(new_n472), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(G15gat), .B1(new_n629), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n475), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(G15gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n629), .B2(new_n644), .ZN(G1326gat));
  NAND2_X1  g444(.A1(new_n632), .A2(new_n437), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT99), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  INV_X1    g448(.A(new_n627), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n543), .A2(new_n574), .A3(new_n606), .A4(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n651), .A2(G29gat), .A3(new_n430), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT45), .Z(new_n653));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n410), .A2(new_n426), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n414), .B(new_n423), .C1(new_n655), .C2(new_n425), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n403), .A2(new_n391), .A3(new_n400), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n437), .B1(new_n657), .B2(new_n345), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n656), .A2(new_n658), .B1(new_n436), .B2(new_n437), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n481), .B1(new_n659), .B2(new_n641), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n660), .B2(new_n605), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n605), .A2(new_n654), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n474), .B2(new_n481), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n574), .A2(new_n541), .A3(new_n650), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT100), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G29gat), .B1(new_n666), .B2(new_n430), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n653), .A2(new_n667), .ZN(G1328gat));
  INV_X1    g467(.A(new_n345), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n651), .A2(G36gat), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT46), .ZN(new_n671));
  OAI21_X1  g470(.A(G36gat), .B1(new_n666), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1329gat));
  OAI21_X1  g472(.A(G43gat), .B1(new_n666), .B2(new_n641), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n643), .A2(G43gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n651), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g476(.A1(new_n651), .A2(new_n265), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n437), .A2(G50gat), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n678), .A2(G50gat), .B1(new_n666), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g480(.A(new_n574), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n542), .A3(new_n605), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n650), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT101), .Z(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n660), .ZN(new_n686));
  INV_X1    g485(.A(new_n430), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(new_n544), .Z(G1332gat));
  AOI21_X1  g488(.A(new_n669), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT102), .Z(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1333gat));
  OAI21_X1  g493(.A(new_n686), .B1(new_n639), .B2(new_n640), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n643), .A2(G71gat), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n695), .A2(G71gat), .B1(new_n686), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g497(.A1(new_n686), .A2(new_n437), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G78gat), .ZN(G1335gat));
  OR3_X1    g499(.A1(new_n682), .A2(KEYINPUT103), .A3(new_n541), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT103), .B1(new_n682), .B2(new_n541), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n650), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n473), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n467), .A2(new_n472), .A3(KEYINPUT98), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n428), .A2(new_n705), .A3(new_n438), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n477), .A2(new_n480), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n605), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n663), .B(new_n703), .C1(new_n711), .C2(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n661), .A2(KEYINPUT104), .A3(new_n663), .A4(new_n703), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716), .B2(new_n430), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n710), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n606), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n701), .A2(new_n702), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT51), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n627), .A2(new_n576), .A3(new_n687), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(G1336gat));
  NOR3_X1   g524(.A1(new_n650), .A2(new_n669), .A3(G92gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n712), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n345), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n712), .B2(new_n669), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n729), .A2(G92gat), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n727), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n714), .A2(new_n345), .A3(new_n715), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n722), .A2(new_n726), .B1(new_n735), .B2(G92gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n716), .B2(new_n641), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n643), .A2(G99gat), .A3(new_n650), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n723), .B2(new_n741), .ZN(G1338gat));
  NOR3_X1   g541(.A1(new_n650), .A2(new_n265), .A3(G106gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n722), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745));
  OAI21_X1  g544(.A(G106gat), .B1(new_n712), .B2(new_n265), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n714), .A2(new_n437), .A3(new_n715), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G106gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(KEYINPUT107), .B1(new_n722), .B2(new_n743), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n752), .A3(G106gat), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n748), .B(new_n745), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n753), .A3(new_n744), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT108), .B1(new_n756), .B2(KEYINPUT53), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n747), .B1(new_n754), .B2(new_n757), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n534), .A2(new_n535), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n529), .B1(new_n522), .B2(new_n528), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n486), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n540), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n627), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n591), .A2(new_n613), .A3(new_n562), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n615), .A2(new_n617), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n619), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n623), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(new_n619), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n770), .B(KEYINPUT54), .C1(new_n618), .C2(new_n611), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n771), .A3(KEYINPUT55), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n536), .A2(new_n488), .A3(new_n537), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n626), .B(new_n772), .C1(new_n773), .C2(new_n538), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT55), .B1(new_n769), .B2(new_n771), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n764), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n605), .ZN(new_n777));
  INV_X1    g576(.A(new_n775), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n772), .A2(new_n626), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n606), .A2(new_n763), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n682), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n683), .A2(new_n627), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n759), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n541), .A2(new_n778), .A3(new_n779), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n606), .B1(new_n784), .B2(new_n764), .ZN(new_n785));
  AND4_X1   g584(.A1(new_n606), .A2(new_n779), .A3(new_n763), .A4(new_n778), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n574), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n683), .A2(new_n627), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n477), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n345), .A2(new_n430), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n542), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(new_n350), .ZN(G1340gat));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n650), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n348), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT111), .B(G120gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n797), .B2(new_n800), .ZN(G1341gat));
  NOR2_X1   g600(.A1(new_n794), .A2(new_n574), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(G127gat), .Z(G1342gat));
  NOR4_X1   g602(.A1(new_n605), .A2(G134gat), .A3(new_n430), .A4(new_n345), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT112), .Z(new_n806));
  OR2_X1    g605(.A1(new_n806), .A2(KEYINPUT56), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(KEYINPUT56), .ZN(new_n808));
  OAI21_X1  g607(.A(G134gat), .B1(new_n794), .B2(new_n605), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(G1343gat));
  XNOR2_X1  g609(.A(new_n775), .B(KEYINPUT113), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n764), .B1(new_n811), .B2(new_n774), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT114), .B(new_n764), .C1(new_n811), .C2(new_n774), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n605), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n682), .B1(new_n816), .B2(new_n780), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n782), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT57), .B1(new_n818), .B2(new_n265), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n783), .A2(new_n789), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n437), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n641), .A2(new_n793), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n819), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT117), .B1(new_n825), .B2(new_n542), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n815), .A2(new_n605), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n786), .B1(new_n827), .B2(new_n814), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n788), .B1(new_n828), .B2(new_n682), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n437), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(new_n830), .B2(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n541), .A4(new_n822), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n826), .A2(new_n833), .A3(G141gat), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n641), .A2(new_n437), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n687), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(KEYINPUT116), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n790), .A2(KEYINPUT116), .A3(new_n430), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n542), .A2(G141gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n669), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n834), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n841), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n831), .A2(new_n845), .A3(new_n822), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n846), .A3(new_n541), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n843), .B1(new_n847), .B2(G141gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n842), .B1(new_n848), .B2(new_n835), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n838), .A2(new_n839), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n345), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n207), .A3(new_n627), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n844), .A2(new_n846), .A3(new_n627), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n207), .A2(KEYINPUT59), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n817), .B2(new_n782), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n788), .C1(new_n828), .C2(new_n682), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n265), .A2(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n790), .B2(new_n265), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n627), .A3(new_n824), .A4(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT119), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n207), .B1(new_n863), .B2(KEYINPUT119), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n852), .B1(new_n855), .B2(new_n866), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n844), .A2(new_n846), .ZN(new_n868));
  OAI21_X1  g667(.A(G155gat), .B1(new_n868), .B2(new_n574), .ZN(new_n869));
  INV_X1    g668(.A(G155gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n870), .A3(new_n682), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n868), .B2(new_n605), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n605), .A2(G162gat), .A3(new_n345), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n850), .B2(new_n874), .ZN(G1347gat));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n783), .A2(new_n430), .A3(new_n789), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n791), .A2(new_n669), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n541), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G169gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n877), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n783), .A2(new_n789), .A3(KEYINPUT120), .A4(new_n430), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(new_n878), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT121), .B(new_n879), .C1(new_n887), .C2(new_n888), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n541), .A2(new_n279), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n876), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n882), .B(KEYINPUT122), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n889), .A2(new_n878), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n889), .A2(new_n885), .A3(new_n878), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n279), .A3(new_n541), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n894), .A2(new_n900), .ZN(G1348gat));
  NOR4_X1   g700(.A1(new_n877), .A2(new_n280), .A3(new_n650), .A4(new_n879), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n890), .A2(new_n891), .A3(new_n650), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(G176gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n897), .A2(new_n627), .A3(new_n898), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(KEYINPUT124), .A3(new_n280), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n902), .B1(new_n905), .B2(new_n907), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n896), .A2(new_n299), .A3(new_n574), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n295), .B1(new_n880), .B2(new_n682), .ZN(new_n910));
  OR3_X1    g709(.A1(new_n909), .A2(KEYINPUT60), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT60), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1350gat));
  INV_X1    g712(.A(G190gat), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n880), .B2(new_n606), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT61), .Z(new_n916));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n914), .A3(new_n606), .A4(new_n898), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  AND2_X1   g717(.A1(new_n861), .A2(new_n862), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n641), .A2(new_n430), .A3(new_n345), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT126), .Z(new_n921));
  AND2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n542), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n836), .A2(new_n669), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT125), .Z(new_n926));
  NAND3_X1  g725(.A1(new_n889), .A2(new_n541), .A3(new_n926), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n922), .A2(new_n924), .B1(new_n923), .B2(new_n927), .ZN(G1352gat));
  NAND3_X1  g727(.A1(new_n919), .A2(new_n627), .A3(new_n921), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G204gat), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n650), .A2(G204gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n889), .A2(new_n926), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  NOR2_X1   g734(.A1(new_n574), .A2(G211gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n889), .A2(new_n926), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n682), .A3(new_n921), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n606), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G218gat), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n605), .A2(G218gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n889), .A2(new_n926), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1355gat));
endmodule


