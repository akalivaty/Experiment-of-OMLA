

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(KEYINPUT41), .B(n470), .ZN(n484) );
  XNOR2_X1 U327 ( .A(n391), .B(KEYINPUT103), .ZN(n396) );
  XNOR2_X1 U328 ( .A(n306), .B(n305), .ZN(n310) );
  OR2_X1 U329 ( .A1(n392), .A2(n576), .ZN(n368) );
  XNOR2_X1 U330 ( .A(n453), .B(KEYINPUT33), .ZN(n454) );
  INV_X1 U331 ( .A(n439), .ZN(n297) );
  XNOR2_X1 U332 ( .A(n455), .B(n454), .ZN(n457) );
  INV_X1 U333 ( .A(KEYINPUT37), .ZN(n420) );
  XNOR2_X1 U334 ( .A(n298), .B(n297), .ZN(n306) );
  XNOR2_X1 U335 ( .A(n421), .B(n420), .ZN(n528) );
  XOR2_X1 U336 ( .A(n459), .B(n458), .Z(n583) );
  INV_X1 U337 ( .A(G43GAT), .ZN(n461) );
  XNOR2_X1 U338 ( .A(n314), .B(n362), .ZN(n543) );
  XNOR2_X1 U339 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U340 ( .A(n461), .B(KEYINPUT40), .ZN(n462) );
  XNOR2_X1 U341 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n463), .B(n462), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n295) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U346 ( .A(KEYINPUT89), .B(n296), .ZN(n298) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G134GAT), .Z(n300) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT90), .B(G176GAT), .Z(n302) );
  XNOR2_X1 U352 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U354 ( .A(n304), .B(n303), .Z(n305) );
  XOR2_X1 U355 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n308) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT84), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n379) );
  XOR2_X1 U358 ( .A(G15GAT), .B(G127GAT), .Z(n315) );
  XNOR2_X1 U359 ( .A(n379), .B(n315), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U364 ( .A(G169GAT), .B(n313), .ZN(n362) );
  XOR2_X1 U365 ( .A(G8GAT), .B(G183GAT), .Z(n357) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G155GAT), .Z(n347) );
  XOR2_X1 U367 ( .A(n357), .B(n347), .Z(n317) );
  XOR2_X1 U368 ( .A(G1GAT), .B(KEYINPUT71), .Z(n425) );
  XNOR2_X1 U369 ( .A(n425), .B(n315), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n322) );
  XNOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n318) );
  XOR2_X1 U372 ( .A(n318), .B(KEYINPUT72), .Z(n458) );
  XNOR2_X1 U373 ( .A(n458), .B(KEYINPUT83), .ZN(n320) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U376 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U377 ( .A(G64GAT), .B(G78GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U380 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n326) );
  XNOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n492) );
  INV_X1 U385 ( .A(n492), .ZN(n587) );
  XOR2_X1 U386 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n366) );
  XOR2_X1 U387 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n332) );
  XNOR2_X1 U388 ( .A(G218GAT), .B(G106GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U390 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n334) );
  XNOR2_X1 U391 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U393 ( .A(n336), .B(n335), .Z(n346) );
  XNOR2_X1 U394 ( .A(G211GAT), .B(KEYINPUT93), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n337), .B(KEYINPUT92), .ZN(n338) );
  XOR2_X1 U396 ( .A(n338), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U397 ( .A(G197GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n359) );
  XNOR2_X1 U399 ( .A(G78GAT), .B(KEYINPUT75), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n341), .B(G148GAT), .ZN(n456) );
  XOR2_X1 U401 ( .A(KEYINPUT22), .B(n456), .Z(n343) );
  NAND2_X1 U402 ( .A1(G228GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n359), .B(n344), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U406 ( .A(n348), .B(n347), .Z(n352) );
  XOR2_X1 U407 ( .A(G50GAT), .B(G162GAT), .Z(n403) );
  XOR2_X1 U408 ( .A(KEYINPUT2), .B(KEYINPUT94), .Z(n350) );
  XNOR2_X1 U409 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n383) );
  XNOR2_X1 U411 ( .A(n403), .B(n383), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n478) );
  XOR2_X1 U413 ( .A(G92GAT), .B(G218GAT), .Z(n354) );
  XNOR2_X1 U414 ( .A(G36GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n414) );
  XOR2_X1 U416 ( .A(KEYINPUT99), .B(n414), .Z(n356) );
  NAND2_X1 U417 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n358) );
  XOR2_X1 U419 ( .A(n358), .B(n357), .Z(n361) );
  XOR2_X2 U420 ( .A(G176GAT), .B(G64GAT), .Z(n438) );
  XNOR2_X1 U421 ( .A(n359), .B(n438), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n531) );
  NOR2_X1 U424 ( .A1(n543), .A2(n531), .ZN(n364) );
  NOR2_X1 U425 ( .A1(n478), .A2(n364), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n531), .B(KEYINPUT27), .ZN(n392) );
  NAND2_X1 U428 ( .A1(n478), .A2(n543), .ZN(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT26), .B(n367), .ZN(n576) );
  NAND2_X1 U430 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n370), .B(KEYINPUT102), .ZN(n390) );
  XOR2_X1 U432 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n372) );
  XNOR2_X1 U433 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n389) );
  XOR2_X1 U435 ( .A(G155GAT), .B(G120GAT), .Z(n374) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(G127GAT), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U438 ( .A(G85GAT), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(G29GAT), .B(G148GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n387) );
  XOR2_X1 U442 ( .A(G134GAT), .B(KEYINPUT80), .Z(n410) );
  XOR2_X1 U443 ( .A(n410), .B(n379), .Z(n381) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n382), .B(G57GAT), .Z(n385) );
  XNOR2_X1 U447 ( .A(n383), .B(KEYINPUT98), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n573) );
  NAND2_X1 U451 ( .A1(n390), .A2(n573), .ZN(n391) );
  NOR2_X1 U452 ( .A1(n573), .A2(n392), .ZN(n393) );
  XOR2_X1 U453 ( .A(KEYINPUT100), .B(n393), .Z(n540) );
  XOR2_X1 U454 ( .A(n478), .B(KEYINPUT28), .Z(n541) );
  NAND2_X1 U455 ( .A1(n541), .A2(n543), .ZN(n394) );
  NOR2_X1 U456 ( .A1(n540), .A2(n394), .ZN(n395) );
  NOR2_X1 U457 ( .A1(n396), .A2(n395), .ZN(n494) );
  NOR2_X1 U458 ( .A1(n587), .A2(n494), .ZN(n419) );
  XNOR2_X1 U459 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n397), .B(G29GAT), .ZN(n398) );
  XOR2_X1 U461 ( .A(n398), .B(KEYINPUT70), .Z(n400) );
  XNOR2_X1 U462 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n435) );
  XOR2_X1 U464 ( .A(KEYINPUT76), .B(G85GAT), .Z(n402) );
  XNOR2_X1 U465 ( .A(G99GAT), .B(G106GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n452) );
  XOR2_X1 U467 ( .A(n452), .B(n403), .Z(n405) );
  NAND2_X1 U468 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n435), .B(n406), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT79), .B(KEYINPUT64), .Z(n408) );
  XNOR2_X1 U472 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U474 ( .A(n409), .B(KEYINPUT67), .Z(n412) );
  XNOR2_X1 U475 ( .A(n410), .B(KEYINPUT65), .ZN(n411) );
  XNOR2_X1 U476 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U477 ( .A(n413), .B(KEYINPUT9), .Z(n416) );
  XNOR2_X1 U478 ( .A(n414), .B(KEYINPUT10), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n567) );
  XNOR2_X1 U481 ( .A(KEYINPUT81), .B(n567), .ZN(n552) );
  XNOR2_X1 U482 ( .A(KEYINPUT36), .B(n552), .ZN(n589) );
  NAND2_X1 U483 ( .A1(n419), .A2(n589), .ZN(n421) );
  XOR2_X1 U484 ( .A(G141GAT), .B(G197GAT), .Z(n423) );
  XNOR2_X1 U485 ( .A(G36GAT), .B(G50GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n429) );
  XNOR2_X1 U491 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U494 ( .A(G15GAT), .B(G113GAT), .Z(n433) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G22GAT), .ZN(n432) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U498 ( .A(n437), .B(n436), .Z(n513) );
  INV_X1 U499 ( .A(n513), .ZN(n577) );
  XOR2_X1 U500 ( .A(G92GAT), .B(n438), .Z(n441) );
  XNOR2_X1 U501 ( .A(n439), .B(G204GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U503 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n443) );
  XNOR2_X1 U504 ( .A(KEYINPUT31), .B(KEYINPUT74), .ZN(n442) );
  XOR2_X1 U505 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n449) );
  INV_X1 U507 ( .A(n449), .ZN(n447) );
  NAND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n448) );
  INV_X1 U509 ( .A(n448), .ZN(n446) );
  NAND2_X1 U510 ( .A1(n447), .A2(n446), .ZN(n451) );
  NAND2_X1 U511 ( .A1(n449), .A2(n448), .ZN(n450) );
  NAND2_X1 U512 ( .A1(n451), .A2(n450), .ZN(n455) );
  XOR2_X1 U513 ( .A(n452), .B(KEYINPUT77), .Z(n453) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n459) );
  INV_X1 U515 ( .A(n583), .ZN(n470) );
  NAND2_X1 U516 ( .A1(n577), .A2(n470), .ZN(n497) );
  NOR2_X1 U517 ( .A1(n528), .A2(n497), .ZN(n460) );
  XOR2_X1 U518 ( .A(KEYINPUT38), .B(n460), .Z(n511) );
  NOR2_X1 U519 ( .A1(n543), .A2(n511), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n577), .A2(n484), .ZN(n464) );
  XNOR2_X1 U521 ( .A(KEYINPUT46), .B(n464), .ZN(n466) );
  AND2_X1 U522 ( .A1(n567), .A2(n492), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT47), .ZN(n474) );
  NAND2_X1 U525 ( .A1(n587), .A2(n589), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n472), .A2(n577), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT48), .B(n475), .ZN(n539) );
  XOR2_X1 U532 ( .A(KEYINPUT121), .B(n531), .Z(n476) );
  NOR2_X1 U533 ( .A1(n539), .A2(n476), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT54), .ZN(n574) );
  INV_X1 U535 ( .A(n478), .ZN(n479) );
  AND2_X1 U536 ( .A1(n573), .A2(n479), .ZN(n480) );
  AND2_X1 U537 ( .A1(n574), .A2(n480), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NOR2_X1 U539 ( .A1(n543), .A2(n482), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT122), .B(n483), .ZN(n571) );
  NAND2_X1 U541 ( .A1(n571), .A2(n484), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n485) );
  XNOR2_X1 U543 ( .A(n485), .B(G176GAT), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1349GAT) );
  NAND2_X1 U545 ( .A1(n571), .A2(n552), .ZN(n491) );
  XOR2_X1 U546 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n489) );
  XNOR2_X1 U547 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n488) );
  NOR2_X1 U548 ( .A1(n552), .A2(n492), .ZN(n493) );
  XNOR2_X1 U549 ( .A(n493), .B(KEYINPUT16), .ZN(n496) );
  INV_X1 U550 ( .A(n494), .ZN(n495) );
  NAND2_X1 U551 ( .A1(n496), .A2(n495), .ZN(n514) );
  OR2_X1 U552 ( .A1(n497), .A2(n514), .ZN(n505) );
  NOR2_X1 U553 ( .A1(n573), .A2(n505), .ZN(n499) );
  XNOR2_X1 U554 ( .A(KEYINPUT104), .B(KEYINPUT34), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n500), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n531), .A2(n505), .ZN(n502) );
  XNOR2_X1 U558 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n502), .B(n501), .ZN(G1325GAT) );
  NOR2_X1 U560 ( .A1(n543), .A2(n505), .ZN(n504) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  NOR2_X1 U563 ( .A1(n541), .A2(n505), .ZN(n506) );
  XOR2_X1 U564 ( .A(G22GAT), .B(n506), .Z(G1327GAT) );
  NOR2_X1 U565 ( .A1(n511), .A2(n573), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n507), .B(KEYINPUT39), .ZN(n508) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(n508), .ZN(G1328GAT) );
  NOR2_X1 U568 ( .A1(n531), .A2(n511), .ZN(n509) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n509), .Z(n510) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n510), .ZN(G1329GAT) );
  NOR2_X1 U571 ( .A1(n541), .A2(n511), .ZN(n512) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NAND2_X1 U573 ( .A1(n484), .A2(n513), .ZN(n527) );
  NOR2_X1 U574 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U575 ( .A(n515), .B(KEYINPUT107), .ZN(n523) );
  NOR2_X1 U576 ( .A1(n573), .A2(n523), .ZN(n517) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U579 ( .A(G57GAT), .B(n518), .Z(G1332GAT) );
  NOR2_X1 U580 ( .A1(n531), .A2(n523), .ZN(n520) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NOR2_X1 U583 ( .A1(n543), .A2(n523), .ZN(n521) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n541), .A2(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n526), .Z(G1335GAT) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(n529), .Z(n536) );
  NOR2_X1 U592 ( .A1(n536), .A2(n573), .ZN(n530) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  XNOR2_X1 U594 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n531), .A2(n536), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U597 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n543), .A2(n536), .ZN(n535) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n535), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n541), .A2(n536), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n537), .Z(n538) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n557) );
  NAND2_X1 U604 ( .A1(n541), .A2(n557), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT115), .B(n544), .Z(n553) );
  NAND2_X1 U607 ( .A1(n553), .A2(n577), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n545), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n547) );
  NAND2_X1 U610 ( .A1(n553), .A2(n484), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G120GAT), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n550) );
  NAND2_X1 U614 ( .A1(n553), .A2(n587), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n556), .ZN(G1343GAT) );
  INV_X1 U621 ( .A(n576), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U623 ( .A(n559), .B(KEYINPUT119), .Z(n566) );
  INV_X1 U624 ( .A(n566), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n577), .A2(n564), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U628 ( .A1(n564), .A2(n484), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n587), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT120), .B(n568), .Z(n569) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n571), .A2(n587), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n590) );
  NAND2_X1 U643 ( .A1(n590), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n580), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n590), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NAND2_X1 U652 ( .A1(n590), .A2(n587), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

