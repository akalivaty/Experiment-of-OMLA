//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G200), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT67), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n247));
  AND2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G107), .ZN(new_n251));
  INV_X1    g0051(.A(G238), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(G1698), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n249), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT66), .A2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT66), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n257), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(G244), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n243), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n259), .A2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n259), .A2(KEYINPUT70), .A3(G190), .A4(new_n270), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n215), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G77), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n279), .A2(new_n281), .B1(G77), .B2(new_n277), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT15), .B(G87), .Z(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n207), .A3(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT69), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n207), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n284), .B1(new_n207), .B2(new_n285), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n278), .A2(new_n215), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n282), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n276), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G179), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n259), .A2(new_n296), .A3(new_n270), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n294), .B1(new_n273), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n275), .A2(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n263), .A2(new_n265), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n268), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(G223), .B2(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n248), .A2(G222), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n257), .B1(new_n306), .B2(new_n285), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n296), .ZN(new_n312));
  INV_X1    g0112(.A(G150), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n290), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n203), .A2(G20), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT68), .B1(new_n287), .B2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(new_n207), .A3(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n315), .B1(new_n319), .B2(new_n291), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n293), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n279), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n323));
  INV_X1    g0123(.A(new_n277), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n323), .B1(new_n202), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n312), .B(new_n326), .C1(G169), .C2(new_n311), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n311), .A2(G190), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n243), .B2(new_n311), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT71), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT9), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n325), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n325), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT71), .B1(new_n321), .B2(new_n325), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT9), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI211_X1 g0137(.A(KEYINPUT10), .B(new_n329), .C1(new_n334), .C2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT10), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n334), .ZN(new_n340));
  INV_X1    g0140(.A(new_n329), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n300), .B(new_n327), .C1(new_n338), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n288), .A2(new_n289), .ZN(new_n346));
  INV_X1    g0146(.A(G68), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(G50), .B1(G20), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n285), .B2(new_n319), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n293), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT11), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT12), .B1(new_n277), .B2(G68), .ZN(new_n354));
  OR3_X1    g0154(.A1(new_n277), .A2(KEYINPUT12), .A3(G68), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(new_n206), .B2(G20), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n354), .A2(new_n355), .B1(new_n322), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n249), .A2(G232), .A3(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n246), .B(new_n247), .C1(new_n304), .C2(new_n305), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n360), .B(new_n361), .C1(new_n302), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n258), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT13), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n266), .B1(G238), .B2(new_n269), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n359), .B(G169), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n364), .A2(new_n366), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n369), .B1(new_n372), .B2(new_n296), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n359), .B1(new_n372), .B2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n358), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n358), .B1(new_n372), .B2(G200), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n367), .A2(new_n368), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT73), .B1(new_n377), .B2(G190), .ZN(new_n378));
  AND4_X1   g0178(.A1(KEYINPUT73), .A2(new_n370), .A3(G190), .A4(new_n371), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT75), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT74), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n257), .A2(G232), .A3(new_n267), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n301), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n301), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(G226), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  INV_X1    g0189(.A(G223), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n362), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n258), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n298), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n301), .A2(new_n384), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n301), .A2(new_n383), .A3(new_n384), .ZN(new_n396));
  AND4_X1   g0196(.A1(G179), .A2(new_n392), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n382), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G169), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n387), .A2(G179), .A3(new_n392), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT75), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n249), .A2(new_n403), .A3(G20), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n306), .B2(new_n207), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(G58), .B(G68), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n346), .A2(G159), .B1(new_n407), .B2(G20), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n403), .B1(new_n249), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n306), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n347), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n408), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n415), .A3(new_n293), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n291), .B1(new_n206), .B2(G20), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n322), .B1(new_n291), .B2(new_n324), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n398), .A2(new_n402), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n398), .A2(new_n422), .A3(new_n402), .A4(new_n419), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n399), .A2(G190), .ZN(new_n424));
  AOI21_X1  g0224(.A(G200), .B1(new_n387), .B2(new_n392), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n416), .B(new_n418), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n399), .A2(new_n243), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G190), .B2(new_n399), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .A3(new_n416), .A4(new_n418), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n421), .A2(new_n423), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n381), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n340), .A2(new_n341), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT10), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n340), .A2(new_n339), .A3(new_n341), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(KEYINPUT72), .A3(new_n327), .A4(new_n300), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n345), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n345), .A2(new_n433), .A3(new_n438), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n206), .A2(G45), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G250), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n265), .A2(G45), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n258), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G244), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  OAI221_X1 g0249(.A(new_n448), .B1(new_n287), .B2(new_n449), .C1(new_n362), .C2(new_n252), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(new_n258), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n274), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G200), .B2(new_n451), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n279), .B1(new_n206), .B2(G33), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G87), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT81), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT19), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n207), .B1(new_n361), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n459), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G87), .A2(G97), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT79), .B1(new_n461), .B2(new_n251), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT80), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n458), .C1(new_n460), .C2(new_n462), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n207), .B(G68), .C1(new_n304), .C2(new_n305), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n457), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n293), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n283), .A2(new_n277), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n456), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n293), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n470), .B1(new_n463), .B2(KEYINPUT80), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n466), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n479), .A2(KEYINPUT81), .A3(new_n474), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n453), .B(new_n455), .C1(new_n476), .C2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT81), .B1(new_n479), .B2(new_n474), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n456), .A3(new_n475), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n482), .A2(new_n483), .B1(new_n283), .B2(new_n454), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n451), .A2(new_n296), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G169), .B2(new_n451), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n481), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  INV_X1    g0288(.A(new_n262), .ZN(new_n489));
  NOR2_X1   g0289(.A1(KEYINPUT66), .A2(G41), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n206), .B(G45), .C1(new_n488), .C2(G41), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n264), .B1(new_n255), .B2(new_n256), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT78), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n260), .A2(new_n262), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n492), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(KEYINPUT78), .A3(new_n494), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n258), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n497), .A2(new_n500), .B1(new_n501), .B2(G257), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT77), .ZN(new_n503));
  INV_X1    g0303(.A(G244), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n362), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n503), .B(new_n507), .C1(new_n362), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n506), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G190), .B(new_n502), .C1(new_n513), .C2(new_n257), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n251), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n251), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n515), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(G20), .B1(G77), .B2(new_n346), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n477), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n324), .A2(new_n516), .ZN(new_n524));
  INV_X1    g0324(.A(new_n454), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT78), .B1(new_n499), .B2(new_n494), .ZN(new_n528));
  AND4_X1   g0328(.A1(KEYINPUT78), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n491), .A2(new_n493), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n257), .ZN(new_n531));
  INV_X1    g0331(.A(G257), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n506), .A2(new_n508), .A3(new_n512), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n258), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n514), .B(new_n527), .C1(new_n535), .C2(new_n243), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n511), .B1(KEYINPUT4), .B2(new_n505), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n257), .B1(new_n537), .B2(new_n508), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n298), .B1(new_n538), .B2(new_n533), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n523), .A2(new_n526), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n296), .B(new_n502), .C1(new_n513), .C2(new_n257), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n487), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n510), .B(new_n207), .C1(G33), .C2(new_n516), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n293), .C1(new_n207), .C2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT20), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n546), .B(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT83), .B1(new_n362), .B2(new_n532), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n248), .A2(new_n550), .A3(G257), .A4(new_n249), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n249), .A2(G264), .A3(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n306), .A2(G303), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n258), .B1(new_n497), .B2(new_n500), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT5), .B1(new_n260), .B2(new_n262), .ZN(new_n559));
  OAI211_X1 g0359(.A(G270), .B(new_n257), .C1(new_n559), .C2(new_n492), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT82), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n563), .A3(G190), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n497), .A2(new_n500), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n555), .B1(new_n551), .B2(new_n549), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n257), .ZN(new_n567));
  OAI21_X1  g0367(.A(G200), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n277), .A2(G116), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n454), .B2(G116), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n548), .A2(new_n564), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n298), .B1(new_n548), .B2(new_n570), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n567), .B2(new_n562), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n572), .B(KEYINPUT21), .C1(new_n567), .C2(new_n562), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n548), .A2(new_n570), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n558), .A2(new_n563), .A3(G179), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n528), .A2(new_n529), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n246), .A2(G250), .A3(new_n247), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G257), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n306), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(G294), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n287), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n258), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n530), .A2(G264), .A3(new_n257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(G169), .B1(new_n581), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n565), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n592), .B2(new_n296), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n249), .A2(new_n207), .A3(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT22), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT22), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n249), .A2(new_n596), .A3(new_n207), .A4(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n287), .A2(new_n449), .A3(G20), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n207), .B2(G107), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n251), .A2(KEYINPUT23), .A3(G20), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n599), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n293), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT25), .B1(new_n324), .B2(new_n251), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n324), .A2(KEYINPUT25), .A3(new_n251), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n454), .A2(G107), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n593), .A2(KEYINPUT84), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n590), .B(new_n613), .C1(new_n592), .C2(new_n296), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n581), .A2(new_n589), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT85), .B1(new_n615), .B2(G200), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n592), .A2(new_n617), .A3(new_n243), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n274), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n607), .A2(new_n611), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n612), .A2(new_n614), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n443), .A2(new_n544), .A3(new_n580), .A4(new_n623), .ZN(G372));
  NAND2_X1  g0424(.A1(new_n400), .A2(new_n401), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n419), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT18), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n419), .A2(new_n625), .A3(new_n422), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n299), .A2(new_n297), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n380), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n375), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n428), .A2(new_n431), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n437), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n327), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n440), .A2(new_n442), .ZN(new_n639));
  INV_X1    g0439(.A(new_n283), .ZN(new_n640));
  OAI22_X1  g0440(.A1(new_n476), .A2(new_n480), .B1(new_n640), .B2(new_n525), .ZN(new_n641));
  INV_X1    g0441(.A(new_n486), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n481), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT86), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n482), .A2(new_n483), .B1(G87), .B2(new_n454), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n641), .A2(new_n642), .B1(new_n647), .B2(new_n453), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT86), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n487), .B2(new_n542), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n620), .A2(new_n622), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n576), .A2(new_n578), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n621), .A2(new_n593), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n575), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n544), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n643), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n638), .B1(new_n639), .B2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G343), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n577), .ZN(new_n669));
  MUX2_X1   g0469(.A(new_n579), .B(new_n580), .S(new_n669), .Z(new_n670));
  AND2_X1   g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n623), .B1(new_n622), .B2(new_n667), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n298), .B1(new_n591), .B2(new_n565), .ZN(new_n673));
  AND4_X1   g0473(.A1(G179), .A2(new_n565), .A3(new_n588), .A4(new_n587), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT84), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n614), .A3(new_n621), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n672), .B1(new_n676), .B2(new_n667), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n621), .A2(new_n593), .A3(new_n667), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n579), .A2(new_n667), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n623), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n498), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n460), .A2(new_n462), .A3(G116), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n206), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n688), .A2(new_n689), .B1(new_n214), .B2(new_n686), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n689), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(new_n645), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n676), .A2(new_n655), .A3(new_n575), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n536), .A2(new_n542), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n648), .A3(new_n654), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n643), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n667), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n700), .B(new_n667), .C1(new_n653), .C2(new_n659), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n535), .A2(G179), .A3(new_n563), .A4(new_n558), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n448), .B1(new_n287), .B2(new_n449), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n362), .A2(new_n252), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n258), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n447), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n588), .A4(new_n587), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT90), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n704), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT90), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n710), .B(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n567), .A2(new_n296), .A3(new_n562), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n535), .A4(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n615), .A2(G179), .A3(new_n451), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n558), .A2(new_n563), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(new_n718), .C1(new_n538), .C2(new_n533), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n712), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n668), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n544), .A2(new_n580), .A3(new_n623), .A4(new_n667), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n703), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n692), .B1(new_n729), .B2(G1), .ZN(G364));
  AND2_X1   g0530(.A1(new_n207), .A2(G13), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n206), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n686), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n671), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G330), .B2(new_n670), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n215), .B1(G20), .B2(new_n298), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n207), .A2(new_n296), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(G190), .A3(new_n243), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n207), .A2(G179), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n740), .A2(G322), .B1(new_n744), .B2(G329), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n738), .A2(new_n742), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n745), .B(new_n306), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n738), .A2(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n274), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n750), .A2(G326), .B1(new_n752), .B2(G303), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n274), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n207), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n749), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI221_X1 g0558(.A(new_n753), .B1(new_n585), .B2(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n741), .A2(new_n274), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT91), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n748), .B(new_n759), .C1(G283), .C2(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n756), .A2(G68), .B1(new_n752), .B2(G87), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n744), .A2(G159), .ZN(new_n768));
  INV_X1    g0568(.A(new_n750), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n767), .B1(KEYINPUT32), .B2(new_n768), .C1(new_n202), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n755), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(KEYINPUT32), .B1(new_n771), .B2(G97), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n306), .B1(new_n740), .B2(G58), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n285), .C2(new_n747), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n764), .A2(new_n251), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n770), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n737), .B1(new_n766), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n737), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n685), .A2(new_n306), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G355), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G116), .B2(new_n210), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n685), .A2(new_n249), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n261), .B2(new_n214), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n238), .A2(new_n261), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n785), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n777), .B(new_n734), .C1(new_n782), .C2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT92), .Z(new_n792));
  INV_X1    g0592(.A(new_n780), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n670), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n736), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  NOR2_X1   g0596(.A1(new_n737), .A2(new_n778), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n734), .B1(G77), .B2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n739), .A2(new_n585), .B1(new_n743), .B2(new_n746), .ZN(new_n800));
  INV_X1    g0600(.A(new_n747), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n249), .B(new_n800), .C1(G116), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n765), .A2(G87), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n771), .A2(G97), .B1(new_n752), .B2(G107), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G283), .A2(new_n756), .B1(new_n750), .B2(G303), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n740), .A2(G143), .B1(new_n801), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n757), .B2(new_n313), .C1(new_n808), .C2(new_n769), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n765), .A2(G68), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n751), .A2(new_n202), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n249), .B1(new_n743), .B2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n815), .C1(G58), .C2(new_n771), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n811), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n809), .A2(new_n810), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n806), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n799), .B1(new_n819), .B2(new_n737), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n275), .A2(new_n295), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n667), .A2(new_n294), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n630), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n631), .A2(new_n667), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n820), .B1(new_n826), .B2(new_n779), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n300), .A2(new_n667), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n653), .B2(new_n659), .ZN(new_n830));
  INV_X1    g0630(.A(new_n643), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n648), .A2(new_n695), .A3(new_n654), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n657), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n646), .A2(new_n650), .A3(new_n652), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n668), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n835), .B2(new_n826), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(KEYINPUT94), .A3(new_n727), .ZN(new_n837));
  INV_X1    g0637(.A(new_n734), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n727), .C2(new_n836), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT94), .B1(new_n836), .B2(new_n727), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n827), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT95), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  OR2_X1    g0643(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n844), .A2(G116), .A3(new_n216), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n285), .B1(G58), .B2(G68), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n214), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n202), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n206), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n375), .A2(new_n668), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n419), .A2(new_n666), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT97), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n432), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT98), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT98), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n432), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n626), .A2(new_n426), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n857), .A2(new_n426), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n420), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n432), .A2(new_n861), .A3(new_n858), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n861), .B1(new_n432), .B2(new_n858), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT38), .B(new_n869), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n856), .B(KEYINPUT39), .C1(new_n870), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n428), .A2(new_n431), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n419), .B(new_n666), .C1(new_n629), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n626), .A2(new_n857), .A3(new_n426), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n867), .A2(new_n420), .B1(new_n879), .B2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT101), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n876), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n873), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n875), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n876), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n873), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n856), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n855), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n890), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n381), .A2(new_n358), .A3(new_n668), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n668), .A2(new_n358), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n375), .A2(new_n380), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n898));
  INV_X1    g0698(.A(new_n824), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n893), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n629), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n666), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT99), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n897), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n830), .B2(new_n824), .ZN(new_n906));
  AOI211_X1 g0706(.A(KEYINPUT99), .B(new_n903), .C1(new_n906), .C2(new_n890), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n892), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT102), .B1(new_n702), .B2(new_n443), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n443), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n637), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n909), .B(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n884), .A2(new_n873), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n726), .A2(KEYINPUT103), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n723), .A2(new_n724), .A3(new_n917), .A4(new_n725), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n825), .B1(new_n894), .B2(new_n896), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n915), .A2(new_n916), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT40), .B1(new_n889), .B2(new_n873), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n920), .A2(KEYINPUT40), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n923), .A2(new_n639), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n923), .B1(new_n639), .B2(new_n924), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(G330), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n206), .B2(new_n731), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n914), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n853), .B1(new_n929), .B2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n781), .B1(new_n210), .B2(new_n640), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n786), .B2(new_n229), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n747), .A2(new_n202), .B1(new_n743), .B2(new_n808), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n306), .B(new_n934), .C1(G150), .C2(new_n740), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n765), .A2(G77), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n750), .A2(G143), .B1(new_n752), .B2(G58), .ZN(new_n937));
  AOI22_X1  g0737(.A1(G68), .A2(new_n771), .B1(new_n756), .B2(G159), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT108), .B1(new_n752), .B2(G116), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT46), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n585), .B2(new_n757), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n765), .A2(G97), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n249), .B1(new_n744), .B2(G317), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n740), .A2(G303), .B1(new_n801), .B2(G283), .ZN(new_n946));
  AOI22_X1  g0746(.A1(G107), .A2(new_n771), .B1(new_n750), .B2(G311), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n944), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n939), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n838), .B(new_n933), .C1(new_n950), .C2(new_n737), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n647), .A2(new_n667), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n831), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n487), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n954), .B2(new_n793), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n695), .B1(new_n527), .B2(new_n667), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n644), .A2(new_n668), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n679), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n683), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n542), .B1(new_n956), .B2(new_n676), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n960), .A2(KEYINPUT42), .B1(new_n667), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(KEYINPUT42), .B2(new_n960), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT105), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n959), .B(new_n966), .Z(new_n967));
  XOR2_X1   g0767(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n968));
  OR2_X1    g0768(.A1(new_n954), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n683), .A2(new_n680), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n958), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n973));
  XOR2_X1   g0773(.A(new_n972), .B(new_n973), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n958), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT44), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n679), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n683), .B1(new_n677), .B2(new_n682), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n671), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n728), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n686), .B(KEYINPUT41), .Z(new_n982));
  OAI21_X1  g0782(.A(new_n732), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT107), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n970), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n970), .B2(new_n983), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n955), .B1(new_n985), .B2(new_n986), .ZN(G387));
  NAND2_X1  g0787(.A1(new_n980), .A2(new_n733), .ZN(new_n988));
  INV_X1    g0788(.A(new_n737), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n739), .A2(new_n202), .B1(new_n747), .B2(new_n347), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n306), .B(new_n990), .C1(G150), .C2(new_n744), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n283), .A2(new_n771), .B1(new_n750), .B2(G159), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n751), .A2(new_n285), .ZN(new_n993));
  INV_X1    g0793(.A(new_n291), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(new_n756), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n944), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n740), .A2(G317), .B1(new_n801), .B2(G303), .ZN(new_n997));
  INV_X1    g0797(.A(G322), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n757), .B2(new_n746), .C1(new_n998), .C2(new_n769), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n771), .A2(G283), .B1(new_n752), .B2(G294), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT110), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n249), .B1(new_n744), .B2(G326), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n449), .C2(new_n764), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n996), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n989), .B1(new_n1010), .B2(KEYINPUT111), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT111), .B2(new_n1010), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n787), .B1(new_n234), .B2(G45), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n687), .B2(new_n783), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n291), .A2(G50), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT50), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n261), .B1(new_n347), .B2(new_n285), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n687), .B(new_n1017), .C1(new_n1016), .C2(new_n1015), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1014), .A2(new_n1018), .B1(G107), .B2(new_n210), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n838), .B1(new_n1019), .B2(new_n781), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1012), .B(new_n1020), .C1(new_n677), .C2(new_n793), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n729), .A2(new_n980), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n686), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n729), .A2(new_n980), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n988), .B(new_n1021), .C1(new_n1023), .C2(new_n1024), .ZN(G393));
  NAND2_X1  g0825(.A1(new_n958), .A2(new_n780), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n781), .B1(new_n516), .B2(new_n210), .C1(new_n787), .C2(new_n241), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n734), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G317), .A2(new_n750), .B1(new_n740), .B2(G311), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n756), .A2(G303), .ZN(new_n1031));
  INV_X1    g0831(.A(G283), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n449), .B2(new_n755), .C1(new_n1032), .C2(new_n751), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n306), .B1(new_n743), .B2(new_n998), .C1(new_n585), .C2(new_n747), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1030), .A2(new_n1033), .A3(new_n775), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g0837(.A(G159), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n769), .A2(new_n313), .B1(new_n1038), .B2(new_n739), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n751), .A2(new_n347), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n755), .A2(new_n285), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G50), .C2(new_n756), .ZN(new_n1043));
  INV_X1    g0843(.A(G143), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n249), .B1(new_n743), .B2(new_n1044), .C1(new_n291), .C2(new_n747), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1040), .A2(new_n1043), .A3(new_n803), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1037), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1028), .B1(new_n1049), .B2(new_n737), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n978), .A2(new_n733), .B1(new_n1026), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n978), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n686), .B1(new_n1052), .B2(new_n1022), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n978), .B1(new_n729), .B2(new_n980), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G390));
  OAI21_X1  g0857(.A(KEYINPUT39), .B1(new_n870), .B2(new_n874), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT100), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n900), .A2(new_n854), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1059), .A2(new_n886), .A3(new_n875), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n915), .A2(new_n854), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n697), .A2(new_n667), .A3(new_n823), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n824), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n897), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n916), .A2(G330), .A3(new_n918), .A4(new_n919), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n726), .A2(G330), .A3(new_n826), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n905), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1068), .A2(new_n1070), .B1(new_n1061), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n916), .A2(G330), .A3(new_n918), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n639), .A2(new_n1075), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n702), .A2(KEYINPUT102), .A3(new_n443), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n638), .B(new_n1076), .C1(new_n1077), .C2(new_n910), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT114), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n916), .A2(new_n1080), .A3(G330), .A4(new_n918), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n826), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n905), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1072), .A2(new_n1065), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1071), .A2(new_n905), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1069), .A2(new_n1086), .B1(new_n830), .B2(new_n824), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1078), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT115), .B1(new_n1074), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1084), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n826), .A3(new_n1081), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1093), .B2(new_n905), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n913), .B(new_n1076), .C1(new_n1094), .C2(new_n1087), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT115), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1069), .B1(new_n1061), .B2(new_n1067), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1061), .A2(new_n1073), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1095), .B(new_n1096), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n906), .A2(new_n855), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n887), .A2(new_n891), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1067), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1070), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1089), .A2(new_n1104), .A3(new_n1098), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1090), .A2(new_n1100), .A3(new_n686), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT116), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1073), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n733), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n1097), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n732), .B1(new_n1061), .B2(new_n1073), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1104), .A2(KEYINPUT116), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1059), .A2(new_n886), .A3(new_n875), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n779), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n739), .A2(new_n449), .B1(new_n747), .B2(new_n516), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n249), .B(new_n1116), .C1(G294), .C2(new_n744), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1042), .B1(G87), .B2(new_n752), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G107), .A2(new_n756), .B1(new_n750), .B2(G283), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1117), .A2(new_n812), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n249), .B1(new_n739), .B2(new_n814), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G125), .B2(new_n744), .ZN(new_n1122));
  OR3_X1    g0922(.A1(new_n751), .A2(KEYINPUT53), .A3(new_n313), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT117), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n801), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT53), .B1(new_n751), .B2(new_n313), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G128), .A2(new_n750), .B1(new_n756), .B2(G137), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n1038), .B2(new_n755), .C1(new_n202), .C2(new_n764), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1120), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT118), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n989), .B1(new_n1131), .B2(KEYINPUT118), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n734), .B1(new_n994), .B2(new_n798), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1115), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT119), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1139), .B(new_n1136), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1106), .B1(new_n1138), .B2(new_n1140), .ZN(G378));
  AOI21_X1  g0941(.A(new_n838), .B1(new_n202), .B2(new_n797), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n640), .A2(new_n747), .B1(new_n251), .B2(new_n739), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n743), .A2(new_n1032), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1143), .A2(new_n249), .A3(new_n498), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n765), .A2(G58), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n993), .B1(G68), .B2(new_n771), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G97), .A2(new_n756), .B1(new_n750), .B2(G116), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n498), .C2(new_n249), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n739), .A2(new_n1155), .B1(new_n747), .B2(new_n808), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G132), .B2(new_n756), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1125), .A2(new_n752), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G150), .A2(new_n771), .B1(new_n750), .B2(G125), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT121), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n744), .C2(G124), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n764), .B2(new_n1038), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1161), .B2(KEYINPUT59), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1154), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n437), .A2(new_n327), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n666), .B1(new_n335), .B2(new_n336), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT55), .Z(new_n1169));
  OR2_X1    g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1142), .B1(new_n989), .B2(new_n1166), .C1(new_n1175), .C2(new_n779), .ZN(new_n1176));
  INV_X1    g0976(.A(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n923), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1175), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n921), .A2(new_n922), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT40), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n922), .B2(new_n915), .ZN(new_n1182));
  OAI211_X1 g0982(.A(G330), .B(new_n1179), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n909), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n907), .B1(new_n1114), .B2(new_n855), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n904), .A3(new_n1178), .A4(new_n1183), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1176), .B1(new_n1188), .B2(new_n732), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n686), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1185), .A2(new_n1187), .A3(KEYINPUT57), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1078), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1105), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1190), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1078), .B1(new_n1074), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1197), .B2(new_n1188), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1189), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n905), .A2(new_n778), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n734), .B1(G68), .B2(new_n798), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(new_n1203));
  OAI22_X1  g1003(.A1(new_n769), .A2(new_n814), .B1(new_n202), .B2(new_n755), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G159), .B2(new_n752), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1125), .A2(new_n756), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n739), .A2(new_n808), .B1(new_n743), .B2(new_n1155), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n306), .B(new_n1207), .C1(G150), .C2(new_n801), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1146), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n739), .A2(new_n1032), .B1(new_n747), .B2(new_n251), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n249), .B(new_n1210), .C1(G303), .C2(new_n744), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n283), .A2(new_n771), .B1(new_n756), .B2(G116), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n750), .A2(G294), .B1(new_n752), .B2(G97), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1211), .A2(new_n936), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n989), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1203), .A2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1196), .A2(new_n733), .B1(new_n1201), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n982), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1095), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1196), .A2(new_n1192), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(G381));
  OR3_X1    g1021(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1136), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1106), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1199), .A3(new_n1225), .ZN(G407));
  INV_X1    g1026(.A(G213), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(G343), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1199), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(G407), .A2(G213), .A3(new_n1229), .ZN(G409));
  XNOR2_X1  g1030(.A(G393), .B(new_n795), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(G387), .A2(new_n1056), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G387), .A2(new_n1056), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(G387), .A2(new_n1056), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G387), .A2(new_n1056), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1231), .A3(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1199), .A2(G378), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1188), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1185), .A2(new_n1187), .A3(KEYINPUT124), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n733), .A3(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1193), .A2(new_n1218), .A3(new_n1187), .A4(new_n1185), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1176), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1225), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1228), .B1(new_n1240), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1094), .A2(new_n1087), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1249), .B2(new_n1078), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1085), .A2(new_n1078), .A3(new_n1088), .A4(KEYINPUT60), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1095), .A2(new_n1251), .A3(new_n686), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G384), .B(new_n1217), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1217), .B1(new_n1252), .B2(new_n1250), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n842), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1247), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1228), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1256), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1228), .A2(KEYINPUT125), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1255), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(G2897), .A3(new_n1228), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1228), .A2(G2897), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1253), .A2(new_n1255), .A3(new_n1267), .A4(new_n1264), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(KEYINPUT61), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1239), .A2(new_n1257), .A3(new_n1262), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1248), .B2(new_n1269), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1260), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1248), .A2(KEYINPUT62), .A3(new_n1256), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1273), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1278), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT62), .B1(new_n1248), .B2(new_n1256), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1271), .B(new_n1280), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1272), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(KEYINPUT127), .B(new_n1272), .C1(new_n1281), .C2(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G405));
  NAND2_X1  g1090(.A1(G375), .A2(new_n1225), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1240), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(new_n1256), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1273), .ZN(G402));
endmodule


