//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006;
  NOR2_X1   g000(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n205), .A2(G183gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n204), .A2(new_n206), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n209), .A2(G190gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n209), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT66), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n226), .A2(KEYINPUT26), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n226), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n223), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n223), .A2(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(new_n224), .A3(new_n225), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n203), .A2(new_n207), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT24), .A3(new_n222), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n232), .A2(new_n236), .A3(new_n238), .A4(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n230), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G120gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G113gat), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G120gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  INV_X1    g049(.A(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n249), .A2(new_n250), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n254), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G120gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n221), .A2(new_n229), .B1(new_n241), .B2(new_n242), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n255), .A2(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G227gat), .ZN(new_n265));
  INV_X1    g064(.A(G233gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT34), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  AOI221_X4 g067(.A(new_n259), .B1(new_n241), .B2(new_n242), .C1(new_n221), .C2(new_n229), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n262), .B1(new_n230), .B2(new_n243), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT34), .ZN(new_n272));
  INV_X1    g071(.A(new_n267), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n268), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT32), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT67), .B(new_n267), .C1(new_n269), .C2(new_n270), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT33), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  XOR2_X1   g082(.A(G15gat), .B(G43gat), .Z(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n282), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  AOI221_X4 g087(.A(new_n277), .B1(KEYINPUT33), .B2(new_n286), .C1(new_n280), .C2(new_n281), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT31), .B(G50gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G228gat), .A2(G233gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT85), .Z(new_n295));
  XNOR2_X1  g094(.A(G141gat), .B(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n296), .A2(new_n297), .B1(KEYINPUT2), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(KEYINPUT73), .A3(new_n298), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n309));
  AND2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT75), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n298), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n300), .A2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(G155gat), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n306), .A2(new_n313), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT69), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n326), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n335), .A2(new_n325), .A3(new_n327), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT70), .B(KEYINPUT29), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n317), .A2(new_n316), .B1(new_n307), .B2(new_n298), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n342), .A3(new_n314), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n301), .A2(new_n303), .A3(new_n297), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n298), .A2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n296), .A2(new_n297), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n308), .A2(new_n312), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n340), .B(new_n343), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n337), .B1(new_n350), .B2(new_n338), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n295), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT3), .B1(new_n354), .B2(KEYINPUT86), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT29), .B1(new_n334), .B2(new_n336), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n324), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n294), .ZN(new_n360));
  INV_X1    g159(.A(new_n338), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n324), .B2(new_n340), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n362), .B2(new_n337), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n352), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G22gat), .ZN(new_n365));
  INV_X1    g164(.A(G22gat), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n352), .B(new_n366), .C1(new_n359), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n293), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n293), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT84), .B(new_n371), .C1(new_n365), .C2(new_n367), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT67), .B1(new_n264), .B2(new_n267), .ZN(new_n374));
  INV_X1    g173(.A(new_n281), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT32), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n286), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n282), .B1(new_n283), .B2(new_n287), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n381));
  NOR4_X1   g180(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT34), .A4(new_n267), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT68), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n276), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n290), .A2(new_n373), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387));
  OAI211_X1 g186(.A(KEYINPUT71), .B(new_n387), .C1(new_n261), .C2(new_n361), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n389), .B1(new_n244), .B2(new_n338), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n244), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n337), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(G64gat), .B(G92gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  OAI21_X1  g197(.A(new_n387), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n244), .A2(new_n389), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n399), .A2(new_n400), .A3(new_n337), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n395), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n398), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n349), .B1(new_n299), .B2(new_n305), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n314), .A2(new_n318), .A3(new_n315), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT2), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT76), .B(G162gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(G155gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT3), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n259), .A3(new_n350), .ZN(new_n416));
  NAND2_X1  g215(.A1(G225gat), .A2(G233gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n313), .B1(new_n347), .B2(new_n346), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n262), .A3(new_n343), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT4), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n422), .B(KEYINPUT83), .C1(new_n421), .C2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  OR3_X1    g225(.A1(new_n421), .A2(KEYINPUT83), .A3(new_n424), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n419), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n421), .A2(KEYINPUT78), .A3(new_n424), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT78), .B1(new_n421), .B2(new_n424), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n420), .A2(new_n262), .A3(new_n432), .A4(new_n343), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT79), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n324), .A2(new_n435), .A3(new_n432), .A4(new_n262), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n418), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n259), .B1(new_n409), .B2(new_n414), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n421), .ZN(new_n441));
  INV_X1    g240(.A(new_n417), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g242(.A(KEYINPUT80), .B(new_n417), .C1(new_n440), .C2(new_n421), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT5), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n428), .B1(new_n438), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT81), .B(KEYINPUT0), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT82), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n440), .A2(new_n421), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT80), .B1(new_n458), .B2(new_n417), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n439), .A3(new_n442), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n426), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n421), .A2(new_n424), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n421), .A2(KEYINPUT78), .A3(new_n424), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n434), .A4(new_n436), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n419), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(new_n455), .A3(new_n428), .A4(new_n452), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n457), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT72), .B1(new_n405), .B2(new_n398), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472));
  INV_X1    g271(.A(new_n398), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n387), .B1(new_n261), .B2(new_n361), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT71), .B1(new_n261), .B2(new_n387), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n337), .B1(new_n476), .B2(new_n388), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n472), .B(new_n473), .C1(new_n477), .C2(new_n401), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n408), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n202), .B1(new_n386), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n482));
  INV_X1    g281(.A(new_n276), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n379), .B2(new_n380), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n408), .A2(new_n470), .A3(new_n479), .ZN(new_n486));
  INV_X1    g285(.A(new_n202), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n373), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n370), .A2(new_n372), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n480), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT36), .B1(new_n482), .B2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n290), .A2(new_n497), .A3(new_n385), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT37), .B1(new_n477), .B2(new_n401), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT87), .A3(new_n473), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n477), .A2(KEYINPUT37), .A3(new_n401), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT87), .B1(new_n500), .B2(new_n473), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT38), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n398), .A2(KEYINPUT38), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n394), .B1(new_n476), .B2(new_n388), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n399), .A2(new_n400), .A3(new_n394), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT37), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n403), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n470), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n408), .A2(new_n479), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n425), .A2(new_n427), .ZN(new_n516));
  INV_X1    g315(.A(new_n416), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n442), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT39), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n458), .B2(new_n417), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n519), .B(new_n442), .C1(new_n516), .C2(new_n517), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n453), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT40), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT40), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n525), .A3(new_n453), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n446), .A2(new_n452), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n529), .A3(new_n373), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n489), .A2(new_n493), .B1(new_n499), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G43gat), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G50gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT15), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT15), .B1(new_n533), .B2(new_n535), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G29gat), .A2(G36gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT91), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT91), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n538), .A2(new_n550), .A3(new_n547), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n546), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n553), .A2(KEYINPUT89), .A3(new_n536), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT89), .B1(new_n553), .B2(new_n536), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G15gat), .B(G22gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT16), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(G1gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(G1gat), .B2(new_n558), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(G8gat), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n549), .A2(new_n551), .B1(new_n555), .B2(new_n554), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n562), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n564), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT18), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n562), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n565), .B(KEYINPUT13), .Z(new_n574));
  AOI22_X1  g373(.A1(new_n570), .A2(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n570), .B2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n563), .B1(new_n557), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n579), .A2(new_n567), .B1(new_n557), .B2(new_n563), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(new_n565), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT93), .B1(new_n570), .B2(new_n571), .ZN(new_n583));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G197gat), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT11), .B(G169gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT12), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n582), .A2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n531), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  OR2_X1    g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G57gat), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT94), .B1(new_n600), .B2(G64gat), .ZN(new_n601));
  INV_X1    g400(.A(G64gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n601), .B1(G57gat), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n600), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n600), .A2(G64gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(G57gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT9), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n596), .A3(new_n597), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n562), .B1(new_n595), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT96), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n595), .ZN(new_n614));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT95), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n620), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n557), .A2(new_n578), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT8), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  OAI21_X1  g429(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n631), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n625), .A2(new_n567), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n635), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n634), .B(new_n638), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n557), .A2(new_n639), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n645), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n636), .A2(new_n651), .A3(new_n610), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n610), .B1(KEYINPUT98), .B2(new_n634), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n634), .A2(KEYINPUT98), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n605), .A3(new_n609), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n652), .B1(new_n658), .B2(new_n651), .ZN(new_n659));
  INV_X1    g458(.A(G230gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n266), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n650), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT10), .B1(new_n654), .B2(new_n657), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT99), .B(new_n663), .C1(new_n664), .C2(new_n652), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n654), .A2(new_n657), .A3(new_n661), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n662), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n659), .A2(new_n661), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n674), .B2(new_n667), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n676), .A2(KEYINPUT100), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(KEYINPUT100), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n624), .A2(new_n649), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n594), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n470), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  INV_X1    g485(.A(new_n515), .ZN(new_n687));
  OR3_X1    g486(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT101), .B1(new_n682), .B2(new_n687), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(G8gat), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  NAND4_X1  g490(.A1(new_n683), .A2(KEYINPUT42), .A3(new_n515), .A4(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n688), .B2(new_n689), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n690), .B(new_n692), .C1(new_n694), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n496), .A2(new_n498), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n682), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n485), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n682), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n594), .A2(new_n494), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n680), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n624), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n679), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n649), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n594), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n470), .A2(G29gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n709), .A2(KEYINPUT102), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT102), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT45), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n531), .B2(new_n649), .ZN(new_n717));
  INV_X1    g516(.A(new_n649), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n529), .A2(new_n373), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(new_n514), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n492), .B1(new_n481), .B2(new_n488), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n593), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n684), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n540), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n727), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n715), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n709), .A2(G36gat), .A3(new_n687), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n724), .A2(new_n515), .A3(new_n725), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n541), .B2(new_n733), .ZN(G1329gat));
  NAND4_X1  g533(.A1(new_n594), .A2(new_n534), .A3(new_n485), .A4(new_n708), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n696), .A3(new_n723), .A4(new_n725), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT47), .B(new_n735), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(G43gat), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n735), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(KEYINPUT47), .B2(new_n742), .ZN(G1330gat));
  NOR4_X1   g542(.A1(new_n702), .A2(G50gat), .A3(new_n649), .A4(new_n707), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n494), .A3(new_n725), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(G50gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g546(.A1(new_n489), .A2(new_n493), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n499), .A2(new_n530), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n593), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n751), .A2(new_n706), .A3(new_n718), .A4(new_n679), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n470), .ZN(new_n754));
  XOR2_X1   g553(.A(KEYINPUT105), .B(G57gat), .Z(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1332gat));
  INV_X1    g555(.A(new_n753), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n687), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT106), .Z(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1333gat));
  XNOR2_X1  g561(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n757), .A2(new_n765), .A3(new_n485), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT107), .B1(new_n753), .B2(new_n699), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n757), .A2(G71gat), .A3(new_n696), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n764), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n771), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT109), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n772), .A3(new_n763), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n757), .A2(new_n494), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n751), .A2(new_n624), .A3(new_n679), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n724), .A2(new_n684), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G85gat), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n751), .A2(new_n624), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n718), .B(new_n788), .C1(new_n721), .C2(new_n722), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n750), .A2(KEYINPUT51), .A3(new_n718), .A4(new_n788), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n679), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n470), .A2(G85gat), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n786), .A2(new_n787), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n790), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n789), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n679), .A2(new_n687), .A3(G92gat), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n724), .A2(new_n515), .A3(new_n782), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n801), .A2(new_n802), .B1(new_n803), .B2(G92gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(G92gat), .ZN(new_n805));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n794), .A2(G92gat), .A3(new_n687), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n797), .A2(new_n804), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  INV_X1    g608(.A(G99gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n810), .A3(new_n485), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n724), .A2(new_n696), .A3(new_n782), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n810), .ZN(G1338gat));
  NAND4_X1  g612(.A1(new_n717), .A2(new_n494), .A3(new_n723), .A4(new_n782), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n679), .A2(G106gat), .A3(new_n373), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g619(.A(new_n818), .B(new_n820), .C1(new_n791), .C2(new_n792), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n791), .A2(new_n792), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT113), .B1(new_n822), .B2(new_n819), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n817), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n799), .A2(new_n800), .A3(new_n819), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n816), .B1(new_n825), .B2(new_n815), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n815), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  INV_X1    g629(.A(new_n823), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n822), .A2(KEYINPUT113), .A3(new_n819), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n829), .B(new_n830), .C1(new_n833), .C2(new_n817), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n827), .A2(new_n834), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n670), .B1(new_n674), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n662), .A2(KEYINPUT54), .A3(new_n665), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(new_n659), .B2(new_n661), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n664), .A2(KEYINPUT115), .A3(new_n652), .A4(new_n663), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n837), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n662), .A2(new_n665), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n843), .A2(new_n844), .B1(new_n846), .B2(new_n672), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n845), .B(new_n847), .C1(new_n591), .C2(new_n592), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n580), .A2(new_n565), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n573), .A2(new_n574), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n587), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g650(.A(new_n851), .B1(new_n588), .B2(new_n582), .C1(new_n677), .C2(new_n678), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n718), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n845), .A2(new_n847), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n582), .B2(new_n588), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n855), .A3(new_n649), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n706), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n681), .A2(new_n593), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n470), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n386), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n687), .A3(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(G113gat), .A3(new_n593), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n515), .A2(new_n470), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n699), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n857), .A2(new_n858), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT116), .A3(new_n373), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT116), .B1(new_n866), .B2(new_n373), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n751), .B(new_n865), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n870), .B2(G113gat), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT117), .ZN(G1340gat));
  OAI21_X1  g671(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n245), .A3(new_n679), .ZN(new_n874));
  INV_X1    g673(.A(new_n861), .ZN(new_n875));
  INV_X1    g674(.A(new_n679), .ZN(new_n876));
  AOI21_X1  g675(.A(G120gat), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n877), .ZN(G1341gat));
  OAI21_X1  g677(.A(G127gat), .B1(new_n873), .B2(new_n706), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n875), .A2(new_n253), .A3(new_n624), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1342gat));
  OAI21_X1  g680(.A(G134gat), .B1(new_n873), .B2(new_n649), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n718), .A2(new_n687), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT118), .Z(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n859), .A2(new_n251), .A3(new_n860), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n887), .A3(new_n888), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n696), .A2(new_n864), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n373), .B1(new_n857), .B2(new_n858), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n300), .B1(new_n897), .B2(new_n751), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n696), .A2(new_n373), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n859), .A2(new_n687), .A3(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n900), .A2(G141gat), .A3(new_n593), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT58), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n896), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n892), .A2(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n890), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G141gat), .B1(new_n905), .B2(new_n593), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(new_n901), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n909), .ZN(G1344gat));
  OR3_X1    g709(.A1(new_n900), .A2(G148gat), .A3(new_n679), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n680), .B2(new_n751), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n681), .A2(KEYINPUT121), .A3(new_n593), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n857), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n494), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n894), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n892), .A2(new_n919), .A3(KEYINPUT57), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n876), .B1(new_n891), .B2(KEYINPUT119), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(KEYINPUT119), .B2(new_n891), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n912), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT59), .B(new_n302), .C1(new_n897), .C2(new_n876), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n911), .B1(new_n926), .B2(new_n927), .ZN(G1345gat));
  NOR2_X1   g727(.A1(new_n900), .A2(new_n706), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n930));
  AOI21_X1  g729(.A(G155gat), .B1(new_n929), .B2(KEYINPUT122), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n624), .A2(G155gat), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n930), .A2(new_n931), .B1(new_n897), .B2(new_n932), .ZN(G1346gat));
  OAI21_X1  g732(.A(new_n412), .B1(new_n905), .B2(new_n649), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n859), .A2(new_n899), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n884), .A2(new_n412), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(G1347gat));
  AOI21_X1  g736(.A(new_n684), .B1(new_n857), .B2(new_n858), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n386), .A2(new_n687), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n751), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n687), .B2(new_n684), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n515), .A2(new_n944), .A3(new_n470), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n943), .A2(new_n485), .A3(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n866), .A2(new_n373), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT116), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n947), .B1(new_n950), .B2(new_n867), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n593), .A2(new_n224), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(G1348gat));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n225), .A3(new_n876), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n951), .A2(new_n876), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n225), .ZN(G1349gat));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n941), .A2(new_n215), .A3(new_n217), .A4(new_n624), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n951), .A2(new_n624), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n957), .B(new_n958), .C1(new_n959), .C2(new_n203), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n203), .B1(new_n951), .B2(new_n624), .ZN(new_n961));
  INV_X1    g760(.A(new_n958), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT60), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(G1350gat));
  NAND3_X1  g763(.A1(new_n941), .A2(new_n207), .A3(new_n718), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n718), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(G190gat), .ZN(new_n968));
  AOI211_X1 g767(.A(KEYINPUT61), .B(new_n207), .C1(new_n951), .C2(new_n718), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1351gat));
  NAND2_X1  g769(.A1(new_n899), .A2(new_n515), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT124), .Z(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n938), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n751), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n697), .A2(new_n945), .A3(new_n943), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n922), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n751), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  NAND2_X1  g781(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n892), .A2(new_n919), .A3(KEYINPUT57), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n983), .A2(new_n984), .B1(new_n894), .B2(new_n917), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n978), .A2(new_n876), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT126), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n922), .A2(new_n988), .A3(new_n876), .A4(new_n978), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(G204gat), .A3(new_n989), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n973), .A2(G204gat), .A3(new_n679), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1353gat));
  INV_X1    g792(.A(G211gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n974), .A2(new_n994), .A3(new_n624), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n976), .A2(new_n706), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n922), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT63), .ZN(new_n999));
  AOI211_X1 g798(.A(new_n999), .B(new_n994), .C1(new_n922), .C2(new_n996), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n995), .B1(new_n998), .B2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(G218gat), .B1(new_n974), .B2(new_n718), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n718), .A2(G218gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1003), .B1(new_n979), .B2(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n922), .A2(new_n1005), .A3(new_n978), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1004), .B2(new_n1006), .ZN(G1355gat));
endmodule


