//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n585, new_n588, new_n590, new_n591,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n462), .A2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT68), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n475), .B(new_n478), .C1(G136), .C2(new_n463), .ZN(G162));
  INV_X1    g054(.A(G138), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n460), .B2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n481), .B(new_n484), .C1(new_n461), .C2(new_n460), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT69), .A2(G114), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT69), .A2(G114), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n487), .B(G2105), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(KEYINPUT69), .A2(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT69), .A2(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n464), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G102), .ZN(new_n494));
  AOI21_X1  g069(.A(KEYINPUT70), .B1(new_n494), .B2(new_n464), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n490), .B(G2104), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n486), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(new_n502), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(G89), .ZN(new_n514));
  NAND2_X1  g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(G168));
  AOI22_X1  g096(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n504), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n507), .A2(new_n524), .B1(new_n509), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n504), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT71), .B(G81), .Z(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n507), .A2(new_n530), .B1(new_n509), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(G153));
  NAND4_X1  g109(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT72), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND4_X1  g113(.A1(G319), .A2(G483), .A3(G661), .A4(new_n538), .ZN(G188));
  AOI22_X1  g114(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G91), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n504), .B1(new_n541), .B2(new_n507), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT9), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G299));
  INV_X1    g123(.A(G171), .ZN(G301));
  INV_X1    g124(.A(G168), .ZN(G286));
  INV_X1    g125(.A(G166), .ZN(G303));
  OAI21_X1  g126(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n502), .A2(new_n506), .A3(G87), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n506), .A2(G49), .A3(G543), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(G288));
  INV_X1    g130(.A(new_n507), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G86), .ZN(new_n557));
  INV_X1    g132(.A(G61), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n500), .B2(new_n501), .ZN(new_n559));
  AND2_X1   g134(.A1(G73), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n557), .A2(new_n561), .A3(new_n562), .ZN(G305));
  INV_X1    g138(.A(new_n509), .ZN(new_n564));
  AOI22_X1  g139(.A1(G85), .A2(new_n556), .B1(new_n564), .B2(G47), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G290));
  NAND2_X1  g144(.A1(G301), .A2(G868), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(G92), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n507), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT76), .B1(new_n507), .B2(new_n572), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT10), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G54), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n576), .A2(new_n504), .B1(new_n577), .B2(new_n509), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n573), .A2(KEYINPUT10), .A3(new_n574), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n571), .B1(new_n582), .B2(G868), .ZN(G321));
  XOR2_X1   g158(.A(G321), .B(KEYINPUT77), .Z(G284));
  NAND2_X1  g159(.A1(G286), .A2(G868), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n547), .B2(G868), .ZN(G297));
  OAI21_X1  g161(.A(new_n585), .B1(new_n547), .B2(G868), .ZN(G280));
  XNOR2_X1  g162(.A(KEYINPUT78), .B(G559), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n582), .B1(G860), .B2(new_n588), .ZN(G148));
  NAND2_X1  g164(.A1(new_n582), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G868), .B2(new_n533), .ZN(G323));
  XNOR2_X1  g167(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g168(.A(new_n462), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n465), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT13), .ZN(new_n597));
  INV_X1    g172(.A(G2100), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  AOI22_X1  g175(.A1(G123), .A2(new_n473), .B1(new_n463), .B2(G135), .ZN(new_n601));
  NOR3_X1   g176(.A1(new_n464), .A2(KEYINPUT79), .A3(G111), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT79), .B1(new_n464), .B2(G111), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n603), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G2096), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n599), .A2(new_n600), .A3(new_n607), .ZN(G156));
  XNOR2_X1  g183(.A(G2427), .B(G2438), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2430), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT15), .B(G2435), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n612), .A2(KEYINPUT14), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(G2443), .B(G2446), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(G2451), .B(G2454), .Z(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n616), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G1341), .B(G1348), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT81), .Z(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G14), .C1(new_n621), .C2(new_n620), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(G401));
  XOR2_X1   g200(.A(G2072), .B(G2078), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT17), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2067), .B(G2678), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n629), .B2(new_n626), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n630), .B1(KEYINPUT82), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(KEYINPUT82), .B2(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(new_n626), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n635), .A2(new_n631), .A3(new_n628), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT18), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n627), .A2(new_n631), .A3(new_n629), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(new_n606), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(G227));
  XOR2_X1   g217(.A(G1956), .B(G2474), .Z(new_n643));
  XOR2_X1   g218(.A(G1961), .B(G1966), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT84), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT19), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(KEYINPUT84), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n648), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n643), .A2(new_n644), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n645), .A3(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n652), .B(new_n656), .C1(new_n653), .C2(new_n655), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1991), .B(G1996), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1981), .B(G1986), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G229));
  MUX2_X1   g239(.A(G24), .B(G290), .S(G16), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1986), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n463), .A2(G131), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n473), .A2(G119), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n464), .A2(G107), .ZN(new_n670));
  OAI21_X1  g245(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  MUX2_X1   g247(.A(G25), .B(new_n672), .S(G29), .Z(new_n673));
  XOR2_X1   g248(.A(KEYINPUT35), .B(G1991), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n673), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(G288), .A2(KEYINPUT88), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n678));
  NAND4_X1  g253(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  MUX2_X1   g255(.A(G23), .B(new_n680), .S(G16), .Z(new_n681));
  XOR2_X1   g256(.A(KEYINPUT33), .B(G1976), .Z(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G1971), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(G6), .B(G305), .S(G16), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT32), .B(G1981), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  NAND3_X1  g266(.A1(new_n683), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n676), .B1(new_n692), .B2(KEYINPUT34), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n667), .B(new_n693), .C1(KEYINPUT34), .C2(new_n692), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT36), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n473), .A2(G129), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT95), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n465), .A2(G105), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT26), .ZN(new_n700));
  AOI211_X1 g275(.A(new_n698), .B(new_n700), .C1(G141), .C2(new_n463), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n704), .B2(G32), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G34), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G29), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G160), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G2084), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n704), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n704), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT29), .Z(new_n717));
  INV_X1    g292(.A(G2090), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2078), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n498), .A2(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n704), .A2(G27), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n706), .A2(new_n707), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n684), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n684), .ZN(new_n727));
  INV_X1    g302(.A(new_n723), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n725), .A2(new_n727), .B1(new_n728), .B2(G2078), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n714), .A2(new_n719), .A3(new_n724), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n731), .A2(new_n704), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n605), .B2(new_n704), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n684), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n684), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(new_n737), .B2(G1966), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n738), .B1(G1966), .B2(new_n737), .C1(new_n725), .C2(new_n727), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT96), .Z(new_n740));
  NOR2_X1   g315(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n684), .A2(G19), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n533), .B2(new_n684), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G1341), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n704), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n463), .A2(G140), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n473), .A2(G128), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n750));
  OR3_X1    g325(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(new_n704), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n582), .A2(G16), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G4), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT89), .B(G1348), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n744), .B(new_n757), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n759), .A2(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT91), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OR3_X1    g339(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT91), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n704), .A2(G33), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n594), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n767), .A2(KEYINPUT93), .A3(new_n464), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT92), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT25), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT93), .B1(new_n767), .B2(new_n464), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n768), .B(new_n773), .C1(G139), .C2(new_n463), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(new_n704), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n717), .A2(new_n718), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n684), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n547), .B2(new_n684), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n776), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n741), .A2(new_n764), .A3(new_n765), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n695), .A2(new_n783), .ZN(G311));
  INV_X1    g359(.A(G311), .ZN(G150));
  NAND2_X1  g360(.A1(new_n582), .A2(G559), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT38), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n504), .ZN(new_n789));
  INV_X1    g364(.A(G93), .ZN(new_n790));
  INV_X1    g365(.A(G55), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n507), .A2(new_n790), .B1(new_n509), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n533), .B(new_n793), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n787), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT39), .ZN(new_n796));
  INV_X1    g371(.A(G860), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(KEYINPUT39), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n793), .A2(new_n797), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT37), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT97), .Z(G145));
  XNOR2_X1  g378(.A(new_n754), .B(new_n498), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n702), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n774), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n596), .B(new_n672), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n473), .A2(G130), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT98), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n463), .A2(G142), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n464), .A2(G118), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n807), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n806), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT99), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n806), .A2(new_n814), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n605), .B(new_n471), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G162), .Z(new_n819));
  NOR3_X1   g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(KEYINPUT99), .B2(new_n815), .ZN(new_n821));
  INV_X1    g396(.A(G37), .ZN(new_n822));
  INV_X1    g397(.A(new_n815), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n819), .B1(new_n823), .B2(new_n817), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(G395));
  XNOR2_X1  g402(.A(G290), .B(G303), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n680), .B(G305), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT42), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n590), .B(new_n794), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n582), .B(new_n547), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(KEYINPUT41), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(KEYINPUT41), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(new_n837), .B2(new_n832), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n831), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G868), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G868), .B2(new_n793), .ZN(G331));
  XOR2_X1   g416(.A(G331), .B(KEYINPUT101), .Z(G295));
  NOR2_X1   g417(.A1(new_n794), .A2(G301), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n533), .B(new_n793), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(G171), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n843), .A2(new_n845), .A3(G286), .ZN(new_n846));
  OAI21_X1  g421(.A(G286), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n835), .B2(new_n836), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n833), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n830), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT104), .B1(new_n849), .B2(new_n850), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n850), .A2(KEYINPUT104), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n830), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n830), .B1(new_n854), .B2(new_n855), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n822), .A3(new_n856), .ZN(new_n863));
  OAI221_X1 g438(.A(KEYINPUT44), .B1(new_n857), .B2(new_n858), .C1(new_n860), .C2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n856), .A2(new_n822), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n860), .B1(new_n866), .B2(new_n861), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n853), .A2(new_n856), .A3(new_n859), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT105), .B1(new_n863), .B2(new_n860), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(G397));
  INV_X1    g448(.A(G1996), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n703), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n754), .B(new_n756), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n702), .A2(G1996), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n879));
  INV_X1    g454(.A(G1384), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT45), .B1(new_n498), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n882), .A2(new_n879), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n672), .B(new_n675), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(G290), .A2(G1986), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n886), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT48), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n754), .A2(new_n756), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n672), .A2(new_n675), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n888), .A2(new_n891), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n703), .B1(new_n896), .B2(G1996), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n886), .B1(new_n897), .B2(new_n876), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n886), .A2(new_n874), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n896), .ZN(new_n901));
  AOI211_X1 g476(.A(KEYINPUT124), .B(KEYINPUT46), .C1(new_n886), .C2(new_n874), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT123), .ZN(new_n907));
  AND2_X1   g482(.A1(G290), .A2(G1986), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n886), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n888), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n498), .A2(new_n880), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT50), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n498), .A2(KEYINPUT109), .A3(new_n880), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(KEYINPUT50), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n879), .A2(G2084), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n880), .ZN(new_n920));
  INV_X1    g495(.A(new_n879), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(G168), .B(new_n919), .C1(new_n925), .C2(G1966), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(G8), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1966), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n913), .B2(new_n915), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n931), .B2(new_n922), .ZN(new_n932));
  AOI21_X1  g507(.A(G168), .B1(new_n932), .B2(new_n919), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n934), .A2(G8), .A3(new_n926), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n929), .B1(new_n935), .B2(KEYINPUT51), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n879), .B1(new_n881), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n920), .A2(KEYINPUT108), .ZN(new_n940));
  INV_X1    g515(.A(new_n497), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n483), .B2(new_n485), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n496), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n939), .A2(new_n940), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n937), .B1(new_n947), .B2(G2078), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n937), .A2(G2078), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n925), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n916), .A2(new_n921), .A3(new_n917), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT121), .B(G1961), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G171), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n940), .A2(new_n945), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(new_n949), .A3(new_n921), .A4(new_n882), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n948), .A2(G301), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT54), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  NOR2_X1   g535(.A1(G166), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n962));
  OR2_X1    g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(KEYINPUT110), .B2(KEYINPUT55), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n921), .B1(new_n911), .B2(KEYINPUT50), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(new_n718), .B1(new_n947), .B2(new_n687), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n970), .B2(new_n960), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n947), .A2(new_n687), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n916), .A2(new_n718), .A3(new_n921), .A4(new_n917), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(G8), .A3(new_n965), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n913), .A2(new_n915), .A3(new_n921), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n677), .A2(G1976), .A3(new_n679), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT52), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT112), .B(G86), .Z(new_n981));
  OAI211_X1 g556(.A(new_n561), .B(new_n562), .C1(new_n507), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G1981), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n557), .A2(new_n984), .A3(new_n561), .A4(new_n562), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n987), .A3(G1981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n990), .A3(new_n988), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(G8), .A3(new_n993), .A4(new_n976), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n978), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n996), .A2(G8), .A3(new_n976), .A4(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n980), .A2(new_n994), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n971), .A2(new_n975), .A3(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n936), .A2(new_n959), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n546), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n543), .A2(new_n545), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n911), .A2(new_n938), .A3(new_n924), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n946), .A2(new_n1010), .A3(new_n921), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n940), .A2(new_n945), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT56), .B(G2072), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n915), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT109), .B1(new_n498), .B2(new_n880), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n968), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1956), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1009), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1956), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n967), .B2(new_n968), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1009), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(new_n947), .C2(new_n1014), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT61), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT61), .A3(new_n1024), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1016), .A2(new_n1017), .A3(new_n879), .ZN(new_n1032));
  INV_X1    g607(.A(G1348), .ZN(new_n1033));
  AOI221_X4 g608(.A(new_n1031), .B1(new_n1032), .B2(new_n756), .C1(new_n951), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT119), .B(G1996), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1011), .A2(new_n1012), .A3(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT58), .B(G1341), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n533), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(KEYINPUT59), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1034), .A2(new_n581), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n951), .A2(new_n1033), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n976), .A2(G2067), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1031), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1033), .B2(new_n951), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT60), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n582), .A3(new_n1047), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1049));
  OR2_X1    g624(.A1(new_n1039), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1030), .A2(new_n1042), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1023), .B1(new_n947), .B2(new_n1014), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1009), .A2(KEYINPUT117), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1024), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1052), .A2(KEYINPUT118), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n582), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1055), .A2(new_n1053), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT118), .B1(new_n1059), .B2(new_n1052), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1025), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1051), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n948), .A2(new_n953), .A3(new_n957), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G171), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n948), .A2(G301), .A3(new_n950), .A4(new_n953), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT54), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1064), .A2(KEYINPUT122), .A3(KEYINPUT54), .A4(new_n1065), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1002), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n926), .A2(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n933), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n928), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(new_n928), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1001), .A2(new_n955), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(G286), .A2(new_n960), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n932), .B2(new_n919), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n971), .A2(new_n975), .A3(new_n1000), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n975), .A2(new_n1000), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n960), .B1(new_n972), .B2(new_n973), .ZN(new_n1088));
  OAI211_X1 g663(.A(KEYINPUT63), .B(new_n1082), .C1(new_n1088), .C2(new_n965), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n980), .A2(new_n994), .A3(new_n999), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n965), .B2(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n974), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n966), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1082), .A2(KEYINPUT63), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1092), .A2(KEYINPUT115), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1085), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G288), .A2(G1976), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n994), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n985), .ZN(new_n1100));
  INV_X1    g675(.A(new_n977), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n975), .B2(new_n1091), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1079), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n907), .B(new_n910), .C1(new_n1071), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1002), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1076), .B1(new_n1073), .B2(new_n928), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n956), .A2(new_n720), .A3(new_n946), .A4(new_n939), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1110), .A2(new_n937), .B1(new_n951), .B2(new_n952), .ZN(new_n1111));
  AOI21_X1  g686(.A(G301), .B1(new_n1111), .B2(new_n950), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n971), .A3(new_n975), .A4(new_n1000), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1103), .B1(new_n1114), .B2(new_n1077), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1108), .A2(new_n1115), .A3(new_n1097), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n907), .B1(new_n1116), .B2(new_n910), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n906), .B1(new_n1107), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT126), .B(new_n906), .C1(new_n1107), .C2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g697(.A1(G227), .A2(new_n458), .ZN(new_n1124));
  AOI21_X1  g698(.A(KEYINPUT127), .B1(new_n624), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g699(.A1(new_n1125), .A2(G229), .ZN(new_n1126));
  NAND3_X1  g700(.A1(new_n624), .A2(KEYINPUT127), .A3(new_n1124), .ZN(new_n1127));
  AND2_X1   g701(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g702(.A(new_n1128), .B(new_n825), .C1(new_n869), .C2(new_n870), .ZN(G225));
  INV_X1    g703(.A(G225), .ZN(G308));
endmodule


