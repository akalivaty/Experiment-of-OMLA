

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n534), .A2(n533), .ZN(G160) );
  XNOR2_X1 U555 ( .A(KEYINPUT32), .B(KEYINPUT96), .ZN(n666) );
  XNOR2_X1 U556 ( .A(n667), .B(n666), .ZN(n675) );
  NOR2_X2 U557 ( .A1(n594), .A2(n697), .ZN(n639) );
  OR2_X1 U558 ( .A1(KEYINPUT33), .A2(n682), .ZN(n687) );
  NOR2_X1 U559 ( .A1(n583), .A2(n536), .ZN(n774) );
  NOR2_X1 U560 ( .A1(G651), .A2(n583), .ZN(n769) );
  NOR2_X1 U561 ( .A1(n625), .A2(n624), .ZN(n934) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X2 U563 ( .A(KEYINPUT17), .B(n520), .Z(n865) );
  NAND2_X1 U564 ( .A1(G138), .A2(n865), .ZN(n522) );
  INV_X1 U565 ( .A(G2105), .ZN(n523) );
  AND2_X1 U566 ( .A1(n523), .A2(G2104), .ZN(n867) );
  NAND2_X1 U567 ( .A1(G102), .A2(n867), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n523), .ZN(n871) );
  NAND2_X1 U570 ( .A1(G126), .A2(n871), .ZN(n525) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U572 ( .A1(G114), .A2(n872), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U575 ( .A1(n871), .A2(G125), .ZN(n530) );
  NAND2_X1 U576 ( .A1(G101), .A2(n867), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT23), .B(n528), .Z(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U579 ( .A1(G137), .A2(n865), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G113), .A2(n872), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n583) );
  INV_X1 U583 ( .A(G651), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G73), .A2(n774), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT2), .ZN(n544) );
  NOR2_X1 U586 ( .A1(G543), .A2(n536), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n537), .Z(n768) );
  NAND2_X1 U588 ( .A1(G61), .A2(n768), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n773) );
  NAND2_X1 U590 ( .A1(G86), .A2(n773), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G48), .A2(n769), .ZN(n540) );
  XNOR2_X1 U593 ( .A(KEYINPUT77), .B(n540), .ZN(n541) );
  NOR2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n544), .A2(n543), .ZN(G305) );
  NAND2_X1 U596 ( .A1(G64), .A2(n768), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G52), .A2(n769), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n552) );
  NAND2_X1 U599 ( .A1(n774), .A2(G77), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT67), .B(n547), .Z(n549) );
  NAND2_X1 U601 ( .A1(n773), .A2(G90), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U604 ( .A1(n552), .A2(n551), .ZN(G171) );
  INV_X1 U605 ( .A(G171), .ZN(G301) );
  NAND2_X1 U606 ( .A1(G91), .A2(n773), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G78), .A2(n774), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n768), .A2(G65), .ZN(n555) );
  XOR2_X1 U610 ( .A(KEYINPUT68), .B(n555), .Z(n556) );
  NOR2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U612 ( .A1(n769), .A2(G53), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U614 ( .A1(G63), .A2(n768), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G51), .A2(n769), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n562), .ZN(n569) );
  NAND2_X1 U618 ( .A1(n773), .A2(G89), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G76), .A2(n774), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U622 ( .A(KEYINPUT5), .B(n566), .ZN(n567) );
  XNOR2_X1 U623 ( .A(KEYINPUT73), .B(n567), .ZN(n568) );
  NOR2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U625 ( .A(KEYINPUT7), .B(n570), .ZN(n929) );
  XNOR2_X1 U626 ( .A(n929), .B(KEYINPUT8), .ZN(G286) );
  NAND2_X1 U627 ( .A1(G62), .A2(n768), .ZN(n571) );
  XNOR2_X1 U628 ( .A(n571), .B(KEYINPUT78), .ZN(n578) );
  NAND2_X1 U629 ( .A1(G88), .A2(n773), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G75), .A2(n774), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G50), .A2(n769), .ZN(n574) );
  XNOR2_X1 U633 ( .A(KEYINPUT79), .B(n574), .ZN(n575) );
  NOR2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U636 ( .A(KEYINPUT80), .B(n579), .Z(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(G49), .A2(n769), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U641 ( .A1(n768), .A2(n582), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n583), .A2(G87), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n585), .A2(n584), .ZN(G288) );
  NAND2_X1 U644 ( .A1(G60), .A2(n768), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G47), .A2(n769), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U647 ( .A(KEYINPUT66), .B(n588), .ZN(n591) );
  NAND2_X1 U648 ( .A1(G85), .A2(n773), .ZN(n589) );
  XNOR2_X1 U649 ( .A(KEYINPUT65), .B(n589), .ZN(n590) );
  NOR2_X1 U650 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U651 ( .A1(n774), .A2(G72), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n593), .A2(n592), .ZN(G290) );
  NOR2_X1 U653 ( .A1(G164), .A2(G1384), .ZN(n698) );
  INV_X1 U654 ( .A(n698), .ZN(n594) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n697) );
  INV_X1 U656 ( .A(n639), .ZN(n659) );
  NAND2_X1 U657 ( .A1(G8), .A2(n659), .ZN(n691) );
  NOR2_X1 U658 ( .A1(G1981), .A2(G305), .ZN(n595) );
  XOR2_X1 U659 ( .A(n595), .B(KEYINPUT24), .Z(n596) );
  NOR2_X1 U660 ( .A1(n691), .A2(n596), .ZN(n696) );
  NOR2_X1 U661 ( .A1(G1966), .A2(n691), .ZN(n671) );
  NOR2_X1 U662 ( .A1(G2084), .A2(n659), .ZN(n668) );
  NOR2_X1 U663 ( .A1(n671), .A2(n668), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT95), .B(n597), .Z(n598) );
  NAND2_X1 U665 ( .A1(G8), .A2(n598), .ZN(n599) );
  XOR2_X1 U666 ( .A(KEYINPUT30), .B(n599), .Z(n600) );
  NAND2_X1 U667 ( .A1(n600), .A2(n929), .ZN(n604) );
  XOR2_X1 U668 ( .A(G2078), .B(KEYINPUT25), .Z(n908) );
  NOR2_X1 U669 ( .A1(n908), .A2(n659), .ZN(n602) );
  NOR2_X1 U670 ( .A1(n639), .A2(G1961), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n653) );
  NAND2_X1 U672 ( .A1(n653), .A2(G301), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT31), .ZN(n658) );
  NAND2_X1 U675 ( .A1(G79), .A2(n774), .ZN(n612) );
  NAND2_X1 U676 ( .A1(G66), .A2(n768), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G54), .A2(n769), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G92), .A2(n773), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT71), .B(n608), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT15), .ZN(n614) );
  XOR2_X1 U684 ( .A(KEYINPUT72), .B(n614), .Z(n933) );
  NAND2_X1 U685 ( .A1(n659), .A2(G1341), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT92), .ZN(n626) );
  XOR2_X1 U687 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n617) );
  NAND2_X1 U688 ( .A1(G56), .A2(n768), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(n625) );
  NAND2_X1 U690 ( .A1(G68), .A2(n774), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n773), .A2(G81), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT12), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(KEYINPUT13), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G43), .A2(n769), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n626), .A2(n934), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G1996), .A2(n639), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT26), .B(n627), .Z(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT64), .B(n630), .Z(n631) );
  NAND2_X1 U702 ( .A1(n933), .A2(n631), .ZN(n638) );
  OR2_X1 U703 ( .A1(n631), .A2(n933), .ZN(n636) );
  INV_X1 U704 ( .A(G2067), .ZN(n818) );
  NOR2_X1 U705 ( .A1(n659), .A2(n818), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n632), .B(KEYINPUT93), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n659), .A2(G1348), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n645) );
  INV_X1 U711 ( .A(G299), .ZN(n935) );
  NAND2_X1 U712 ( .A1(G1956), .A2(n659), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n639), .A2(G2072), .ZN(n640) );
  XOR2_X1 U714 ( .A(KEYINPUT27), .B(n640), .Z(n641) );
  NAND2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT90), .B(n643), .Z(n646) );
  NAND2_X1 U717 ( .A1(n935), .A2(n646), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n935), .A2(n646), .ZN(n648) );
  XNOR2_X1 U720 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n653), .A2(G301), .ZN(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT89), .B(n654), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n672), .A2(G286), .ZN(n664) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n691), .ZN(n661) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n659), .ZN(n660) );
  NOR2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U733 ( .A1(G303), .A2(n662), .ZN(n663) );
  NAND2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n665), .A2(G8), .ZN(n667) );
  NAND2_X1 U736 ( .A1(G8), .A2(n668), .ZN(n669) );
  XOR2_X1 U737 ( .A(KEYINPUT88), .B(n669), .Z(n670) );
  NOR2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n690) );
  NOR2_X1 U741 ( .A1(G1976), .A2(G288), .ZN(n942) );
  NOR2_X1 U742 ( .A1(G303), .A2(G1971), .ZN(n676) );
  XOR2_X1 U743 ( .A(n676), .B(KEYINPUT97), .Z(n677) );
  NOR2_X1 U744 ( .A1(n942), .A2(n677), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n690), .A2(n678), .ZN(n680) );
  NAND2_X1 U746 ( .A1(G288), .A2(G1976), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n679), .B(KEYINPUT98), .ZN(n943) );
  NAND2_X1 U748 ( .A1(n680), .A2(n943), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n691), .A2(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n942), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n683), .A2(n691), .ZN(n685) );
  XOR2_X1 U752 ( .A(G1981), .B(G305), .Z(n930) );
  INV_X1 U753 ( .A(n930), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n694) );
  NOR2_X1 U756 ( .A1(G2090), .A2(G303), .ZN(n688) );
  NAND2_X1 U757 ( .A1(G8), .A2(n688), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n729) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n743) );
  XOR2_X1 U763 ( .A(KEYINPUT37), .B(n818), .Z(n741) );
  NAND2_X1 U764 ( .A1(G140), .A2(n865), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G104), .A2(n867), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT83), .ZN(n702) );
  XNOR2_X1 U768 ( .A(n702), .B(KEYINPUT34), .ZN(n708) );
  XNOR2_X1 U769 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n706) );
  NAND2_X1 U770 ( .A1(G128), .A2(n871), .ZN(n704) );
  NAND2_X1 U771 ( .A1(G116), .A2(n872), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U773 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U775 ( .A(KEYINPUT36), .B(n709), .Z(n862) );
  NOR2_X1 U776 ( .A1(n741), .A2(n862), .ZN(n998) );
  NAND2_X1 U777 ( .A1(n743), .A2(n998), .ZN(n739) );
  NAND2_X1 U778 ( .A1(G131), .A2(n865), .ZN(n711) );
  NAND2_X1 U779 ( .A1(G95), .A2(n867), .ZN(n710) );
  NAND2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U781 ( .A1(G119), .A2(n871), .ZN(n713) );
  NAND2_X1 U782 ( .A1(G107), .A2(n872), .ZN(n712) );
  NAND2_X1 U783 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n854) );
  XNOR2_X1 U785 ( .A(KEYINPUT85), .B(G1991), .ZN(n903) );
  NOR2_X1 U786 ( .A1(n854), .A2(n903), .ZN(n725) );
  NAND2_X1 U787 ( .A1(G129), .A2(n871), .ZN(n717) );
  NAND2_X1 U788 ( .A1(G117), .A2(n872), .ZN(n716) );
  NAND2_X1 U789 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n867), .A2(G105), .ZN(n718) );
  XOR2_X1 U791 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  NOR2_X1 U792 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U793 ( .A(n721), .B(KEYINPUT86), .ZN(n723) );
  NAND2_X1 U794 ( .A1(G141), .A2(n865), .ZN(n722) );
  NAND2_X1 U795 ( .A1(n723), .A2(n722), .ZN(n861) );
  AND2_X1 U796 ( .A1(n861), .A2(G1996), .ZN(n724) );
  NOR2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n1000) );
  INV_X1 U798 ( .A(n1000), .ZN(n726) );
  NAND2_X1 U799 ( .A1(n726), .A2(n743), .ZN(n733) );
  NAND2_X1 U800 ( .A1(n739), .A2(n733), .ZN(n727) );
  XOR2_X1 U801 ( .A(KEYINPUT87), .B(n727), .Z(n728) );
  NOR2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U803 ( .A(G1986), .B(G290), .ZN(n941) );
  NAND2_X1 U804 ( .A1(n941), .A2(n743), .ZN(n730) );
  NAND2_X1 U805 ( .A1(n731), .A2(n730), .ZN(n746) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n861), .ZN(n732) );
  XOR2_X1 U807 ( .A(KEYINPUT99), .B(n732), .Z(n988) );
  INV_X1 U808 ( .A(n733), .ZN(n736) );
  AND2_X1 U809 ( .A1(n903), .A2(n854), .ZN(n991) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U811 ( .A1(n991), .A2(n734), .ZN(n735) );
  NOR2_X1 U812 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U813 ( .A1(n988), .A2(n737), .ZN(n738) );
  XNOR2_X1 U814 ( .A(n738), .B(KEYINPUT39), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n741), .A2(n862), .ZN(n1002) );
  NAND2_X1 U817 ( .A1(n742), .A2(n1002), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U819 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U820 ( .A(n747), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U821 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U822 ( .A(G57), .ZN(G237) );
  INV_X1 U823 ( .A(G82), .ZN(G220) );
  NAND2_X1 U824 ( .A1(G7), .A2(G661), .ZN(n748) );
  XOR2_X1 U825 ( .A(n748), .B(KEYINPUT10), .Z(n808) );
  NAND2_X1 U826 ( .A1(n808), .A2(G567), .ZN(n749) );
  XOR2_X1 U827 ( .A(KEYINPUT11), .B(n749), .Z(G234) );
  NAND2_X1 U828 ( .A1(n934), .A2(G860), .ZN(G153) );
  INV_X1 U829 ( .A(G868), .ZN(n791) );
  NOR2_X1 U830 ( .A1(G301), .A2(n791), .ZN(n751) );
  NOR2_X1 U831 ( .A1(n933), .A2(G868), .ZN(n750) );
  NOR2_X1 U832 ( .A1(n751), .A2(n750), .ZN(G284) );
  NOR2_X1 U833 ( .A1(G868), .A2(G299), .ZN(n753) );
  NOR2_X1 U834 ( .A1(G286), .A2(n791), .ZN(n752) );
  NOR2_X1 U835 ( .A1(n753), .A2(n752), .ZN(G297) );
  INV_X1 U836 ( .A(G860), .ZN(n780) );
  NAND2_X1 U837 ( .A1(n780), .A2(G559), .ZN(n754) );
  INV_X1 U838 ( .A(n933), .ZN(n881) );
  NAND2_X1 U839 ( .A1(n754), .A2(n881), .ZN(n755) );
  XNOR2_X1 U840 ( .A(n755), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U841 ( .A1(G868), .A2(n881), .ZN(n756) );
  NOR2_X1 U842 ( .A1(G559), .A2(n756), .ZN(n758) );
  AND2_X1 U843 ( .A1(n791), .A2(n934), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(G282) );
  XOR2_X1 U845 ( .A(G2100), .B(KEYINPUT74), .Z(n767) );
  NAND2_X1 U846 ( .A1(G123), .A2(n871), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT18), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n867), .A2(G99), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G135), .A2(n865), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G111), .A2(n872), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n990) );
  XNOR2_X1 U854 ( .A(G2096), .B(n990), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n767), .A2(n766), .ZN(G156) );
  NAND2_X1 U856 ( .A1(G67), .A2(n768), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G55), .A2(n769), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT76), .B(n772), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G93), .A2(n773), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G80), .A2(n774), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n792) );
  NAND2_X1 U864 ( .A1(n881), .A2(G559), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(n934), .ZN(n789) );
  NAND2_X1 U866 ( .A1(n780), .A2(n789), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n781), .B(KEYINPUT75), .ZN(n782) );
  XOR2_X1 U868 ( .A(n792), .B(n782), .Z(G145) );
  XOR2_X1 U869 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n783) );
  XNOR2_X1 U870 ( .A(G288), .B(n783), .ZN(n784) );
  XOR2_X1 U871 ( .A(n792), .B(n784), .Z(n786) );
  XOR2_X1 U872 ( .A(G290), .B(G166), .Z(n785) );
  XNOR2_X1 U873 ( .A(n786), .B(n785), .ZN(n787) );
  XOR2_X1 U874 ( .A(n787), .B(n935), .Z(n788) );
  XNOR2_X1 U875 ( .A(n788), .B(G305), .ZN(n880) );
  XOR2_X1 U876 ( .A(n880), .B(n789), .Z(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n794) );
  NOR2_X1 U878 ( .A1(G868), .A2(n792), .ZN(n793) );
  NOR2_X1 U879 ( .A1(n794), .A2(n793), .ZN(G295) );
  NAND2_X1 U880 ( .A1(G2078), .A2(G2084), .ZN(n796) );
  XOR2_X1 U881 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n795) );
  XNOR2_X1 U882 ( .A(n796), .B(n795), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G2090), .A2(n797), .ZN(n798) );
  XNOR2_X1 U884 ( .A(KEYINPUT21), .B(n798), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n799), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U886 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U887 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U888 ( .A1(G220), .A2(G219), .ZN(n800) );
  XOR2_X1 U889 ( .A(KEYINPUT22), .B(n800), .Z(n801) );
  NOR2_X1 U890 ( .A1(G218), .A2(n801), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G96), .A2(n802), .ZN(n813) );
  NAND2_X1 U892 ( .A1(n813), .A2(G2106), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G69), .A2(G120), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G237), .A2(n803), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G108), .A2(n804), .ZN(n814) );
  NAND2_X1 U896 ( .A1(n814), .A2(G567), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G483), .A2(G661), .ZN(n807) );
  NOR2_X1 U899 ( .A1(n815), .A2(n807), .ZN(n810) );
  NAND2_X1 U900 ( .A1(n810), .A2(G36), .ZN(G176) );
  INV_X1 U901 ( .A(n929), .ZN(G168) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n808), .ZN(G217) );
  INV_X1 U903 ( .A(n808), .ZN(G223) );
  AND2_X1 U904 ( .A1(G15), .A2(G2), .ZN(n809) );
  NAND2_X1 U905 ( .A1(G661), .A2(n809), .ZN(G259) );
  NAND2_X1 U906 ( .A1(G1), .A2(G3), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT100), .ZN(G188) );
  INV_X1 U910 ( .A(G120), .ZN(G236) );
  INV_X1 U911 ( .A(G96), .ZN(G221) );
  INV_X1 U912 ( .A(G69), .ZN(G235) );
  NOR2_X1 U913 ( .A1(n814), .A2(n813), .ZN(G325) );
  INV_X1 U914 ( .A(G325), .ZN(G261) );
  INV_X1 U915 ( .A(n815), .ZN(G319) );
  XOR2_X1 U916 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n817) );
  XNOR2_X1 U917 ( .A(G2678), .B(KEYINPUT43), .ZN(n816) );
  XNOR2_X1 U918 ( .A(n817), .B(n816), .ZN(n822) );
  XOR2_X1 U919 ( .A(KEYINPUT42), .B(G2072), .Z(n820) );
  XOR2_X1 U920 ( .A(n818), .B(G2090), .Z(n819) );
  XNOR2_X1 U921 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U922 ( .A(n822), .B(n821), .Z(n824) );
  XNOR2_X1 U923 ( .A(G2100), .B(G2096), .ZN(n823) );
  XNOR2_X1 U924 ( .A(n824), .B(n823), .ZN(n826) );
  XOR2_X1 U925 ( .A(G2078), .B(G2084), .Z(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(G227) );
  XOR2_X1 U927 ( .A(G1976), .B(G1961), .Z(n828) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1956), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U930 ( .A(G1981), .B(G1966), .Z(n830) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U932 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U933 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U934 ( .A(KEYINPUT103), .B(KEYINPUT41), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n836) );
  XOR2_X1 U936 ( .A(G1971), .B(G2474), .Z(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(G229) );
  NAND2_X1 U938 ( .A1(G124), .A2(n871), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n837), .B(KEYINPUT104), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n838), .B(KEYINPUT44), .ZN(n840) );
  NAND2_X1 U941 ( .A1(G100), .A2(n867), .ZN(n839) );
  NAND2_X1 U942 ( .A1(n840), .A2(n839), .ZN(n844) );
  NAND2_X1 U943 ( .A1(G136), .A2(n865), .ZN(n842) );
  NAND2_X1 U944 ( .A1(G112), .A2(n872), .ZN(n841) );
  NAND2_X1 U945 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U946 ( .A1(n844), .A2(n843), .ZN(G162) );
  NAND2_X1 U947 ( .A1(G130), .A2(n871), .ZN(n846) );
  NAND2_X1 U948 ( .A1(G118), .A2(n872), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G142), .A2(n865), .ZN(n848) );
  NAND2_X1 U951 ( .A1(G106), .A2(n867), .ZN(n847) );
  NAND2_X1 U952 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U953 ( .A(KEYINPUT45), .B(n849), .ZN(n850) );
  XNOR2_X1 U954 ( .A(KEYINPUT105), .B(n850), .ZN(n851) );
  NOR2_X1 U955 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n853), .B(KEYINPUT46), .Z(n856) );
  XNOR2_X1 U957 ( .A(n854), .B(KEYINPUT48), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U959 ( .A(n990), .B(G162), .Z(n858) );
  XNOR2_X1 U960 ( .A(G164), .B(G160), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U963 ( .A(n862), .B(n861), .Z(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n878) );
  NAND2_X1 U965 ( .A1(n865), .A2(G139), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT106), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G103), .A2(n867), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT107), .B(n870), .Z(n877) );
  NAND2_X1 U970 ( .A1(G127), .A2(n871), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n1004) );
  XNOR2_X1 U975 ( .A(n878), .B(n1004), .ZN(n879) );
  NOR2_X1 U976 ( .A1(G37), .A2(n879), .ZN(G395) );
  XOR2_X1 U977 ( .A(G301), .B(n880), .Z(n885) );
  XOR2_X1 U978 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n883) );
  XOR2_X1 U979 ( .A(n881), .B(n934), .Z(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U982 ( .A(G286), .B(n886), .Z(n887) );
  NOR2_X1 U983 ( .A1(G37), .A2(n887), .ZN(G397) );
  XOR2_X1 U984 ( .A(G2451), .B(G2430), .Z(n889) );
  XNOR2_X1 U985 ( .A(G2438), .B(G2443), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n895) );
  XOR2_X1 U987 ( .A(G2435), .B(G2454), .Z(n891) );
  XNOR2_X1 U988 ( .A(G1348), .B(G1341), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n893) );
  XOR2_X1 U990 ( .A(G2446), .B(G2427), .Z(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n896) );
  NAND2_X1 U993 ( .A1(G14), .A2(n896), .ZN(n902) );
  NAND2_X1 U994 ( .A1(G319), .A2(n902), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n897) );
  XNOR2_X1 U996 ( .A(KEYINPUT49), .B(n897), .ZN(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U999 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1000 ( .A(G225), .ZN(G308) );
  INV_X1 U1001 ( .A(G108), .ZN(G238) );
  INV_X1 U1002 ( .A(n902), .ZN(G401) );
  XNOR2_X1 U1003 ( .A(KEYINPUT55), .B(KEYINPUT112), .ZN(n1012) );
  XNOR2_X1 U1004 ( .A(n1012), .B(KEYINPUT118), .ZN(n924) );
  XNOR2_X1 U1005 ( .A(G2090), .B(G35), .ZN(n919) );
  XOR2_X1 U1006 ( .A(G26), .B(G2067), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n903), .B(G25), .ZN(n904) );
  NAND2_X1 U1008 ( .A1(n904), .A2(G28), .ZN(n905) );
  XNOR2_X1 U1009 ( .A(n905), .B(KEYINPUT115), .ZN(n906) );
  NAND2_X1 U1010 ( .A1(n907), .A2(n906), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(G1996), .B(G32), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n908), .B(G27), .ZN(n909) );
  NOR2_X1 U1013 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1014 ( .A(KEYINPUT117), .B(n911), .Z(n914) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(G33), .Z(n912) );
  XNOR2_X1 U1016 ( .A(G2072), .B(n912), .ZN(n913) );
  NAND2_X1 U1017 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1018 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(KEYINPUT53), .B(n917), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n922) );
  XOR2_X1 U1021 ( .A(G2084), .B(KEYINPUT54), .Z(n920) );
  XNOR2_X1 U1022 ( .A(G34), .B(n920), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(G29), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(n926), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n927), .A2(G11), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(KEYINPUT120), .ZN(n986) );
  INV_X1 U1029 ( .A(G16), .ZN(n982) );
  XOR2_X1 U1030 ( .A(n982), .B(KEYINPUT56), .Z(n955) );
  XOR2_X1 U1031 ( .A(n929), .B(G1966), .Z(n931) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(n932), .B(KEYINPUT57), .ZN(n953) );
  XOR2_X1 U1034 ( .A(G1348), .B(n933), .Z(n939) );
  XOR2_X1 U1035 ( .A(n934), .B(G1341), .Z(n937) );
  XOR2_X1 U1036 ( .A(n935), .B(G1956), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n949) );
  INV_X1 U1040 ( .A(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT121), .B(n945), .Z(n947) );
  XOR2_X1 U1043 ( .A(G1971), .B(G166), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1046 ( .A(G1961), .B(G171), .Z(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n984) );
  XNOR2_X1 U1050 ( .A(KEYINPUT123), .B(G1341), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(G19), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT59), .B(G4), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT125), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G1348), .B(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G1956), .B(G20), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT124), .B(G1981), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G6), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT126), .B(n966), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(n967), .B(KEYINPUT60), .ZN(n977) );
  XNOR2_X1 U1063 ( .A(G1961), .B(KEYINPUT122), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(G5), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1971), .B(G22), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(G23), .B(G1976), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1068 ( .A(G1986), .B(G24), .Z(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(KEYINPUT58), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G21), .B(G1966), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT61), .B(n980), .ZN(n981) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n1017) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n989), .Z(n996) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1083 ( .A(KEYINPUT110), .B(n992), .Z(n994) );
  XOR2_X1 U1084 ( .A(G2084), .B(G160), .Z(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT111), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XOR2_X1 U1091 ( .A(G2072), .B(n1004), .Z(n1006) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT50), .B(n1007), .Z(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1010), .Z(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT113), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(n1015), .B(KEYINPUT114), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1018), .ZN(G150) );
  INV_X1 U1103 ( .A(G150), .ZN(G311) );
endmodule

