//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(KEYINPUT67), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT67), .B1(new_n467), .B2(new_n470), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n465), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g053(.A1(new_n472), .A2(new_n473), .A3(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n466), .A2(G136), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n465), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT68), .Z(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n463), .A2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n481), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI211_X1 g067(.A(KEYINPUT70), .B(new_n489), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  XNOR2_X1  g071(.A(new_n496), .B(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n482), .A2(G126), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n492), .B1(new_n499), .B2(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n466), .B(new_n500), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n493), .A2(new_n497), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n506), .A2(new_n507), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n514), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT72), .B1(new_n514), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n505), .B1(KEYINPUT6), .B2(new_n510), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n513), .A2(new_n523), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n515), .A2(new_n518), .ZN(new_n530));
  AND2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(new_n517), .B2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n529), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(new_n519), .A3(KEYINPUT72), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n534), .A2(G89), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(G51), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n536), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n531), .A2(new_n532), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n525), .A2(G52), .B1(new_n547), .B2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n534), .A2(new_n535), .ZN(new_n549));
  INV_X1    g124(.A(G90), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n522), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n545), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n525), .A2(G43), .B1(new_n559), .B2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT78), .ZN(new_n567));
  XOR2_X1   g142(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND3_X1  g145(.A1(new_n519), .A2(G53), .A3(new_n524), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n510), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n534), .A2(G91), .A3(new_n535), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  NAND2_X1  g152(.A1(new_n522), .A2(G87), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n508), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(G49), .A2(new_n525), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n545), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n525), .A2(G48), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n549), .B2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n545), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n525), .A2(G47), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n549), .B2(new_n592), .ZN(G290));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NOR2_X1   g169(.A1(G301), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT79), .B(G66), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n508), .A2(new_n596), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n510), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n525), .A2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT10), .B1(new_n522), .B2(G92), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .A4(new_n535), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n601), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(new_n594), .ZN(G284));
  AOI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(new_n594), .ZN(G321));
  NAND2_X1  g183(.A1(G299), .A2(new_n594), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n594), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n594), .B2(G168), .ZN(G280));
  XNOR2_X1  g186(.A(KEYINPUT81), .B(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(G860), .B2(new_n612), .ZN(G148));
  NAND2_X1  g188(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n490), .A2(new_n469), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n466), .A2(G135), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n482), .A2(G123), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n627));
  INV_X1    g202(.A(G111), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n627), .B2(new_n626), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n622), .A2(new_n623), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT83), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n654), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n652), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n654), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n677), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  OR2_X1    g261(.A1(G5), .A2(G16), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(G301), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G1961), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT97), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT31), .B(G11), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT95), .ZN(new_n694));
  INV_X1    g269(.A(G28), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  AOI21_X1  g271(.A(G29), .B1(new_n695), .B2(KEYINPUT30), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NOR2_X1   g274(.A1(G168), .A2(new_n688), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n688), .B2(G21), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n698), .B1(new_n699), .B2(new_n631), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n702), .B2(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n692), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(KEYINPUT98), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT98), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n692), .A2(new_n707), .A3(new_n704), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n606), .A2(new_n688), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G4), .B2(new_n688), .ZN(new_n710));
  INV_X1    g285(.A(G1348), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n690), .A2(G1961), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n711), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n699), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n490), .A2(G127), .ZN(new_n719));
  NAND2_X1  g294(.A1(G115), .A2(G2104), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n481), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n718), .B(new_n721), .C1(G139), .C2(new_n466), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT92), .Z(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n699), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G2072), .ZN(new_n725));
  NOR2_X1   g300(.A1(G160), .A2(new_n699), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G29), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n724), .B2(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n688), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n562), .B2(new_n688), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NOR2_X1   g311(.A1(G27), .A2(G29), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G164), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n725), .A2(new_n733), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(G29), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n742), .B(new_n746), .C1(G29), .C2(new_n743), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n466), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n482), .A2(G128), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n481), .A2(G116), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n699), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT91), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT91), .ZN(new_n761));
  AOI21_X1  g336(.A(G2067), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n760), .A2(G2067), .A3(new_n761), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n762), .B(new_n763), .C1(new_n731), .C2(new_n730), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n482), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n469), .A2(G105), .ZN(new_n769));
  INV_X1    g344(.A(G141), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n491), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT93), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT94), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(KEYINPUT94), .C1(G29), .C2(G32), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT27), .B(G1996), .Z(new_n777));
  AND3_X1   g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n750), .B(new_n764), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n715), .A2(new_n741), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n688), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT23), .ZN(new_n783));
  INV_X1    g358(.A(G299), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n688), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT99), .ZN(new_n786));
  INV_X1    g361(.A(G1956), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n788), .B(new_n789), .C1(new_n748), .C2(new_n749), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT100), .Z(new_n791));
  NAND4_X1  g366(.A1(new_n706), .A2(new_n708), .A3(new_n781), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n688), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(G288), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n688), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n688), .A2(G22), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n688), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G6), .B(G305), .S(G16), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G1971), .B2(new_n800), .ZN(new_n806));
  OR3_X1    g381(.A1(new_n802), .A2(new_n806), .A3(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n482), .A2(G119), .ZN(new_n808));
  NOR2_X1   g383(.A1(G95), .A2(G2105), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT88), .Z(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(new_n481), .B2(G107), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n466), .A2(KEYINPUT87), .A3(G131), .ZN(new_n812));
  AOI21_X1  g387(.A(KEYINPUT87), .B1(new_n466), .B2(G131), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n808), .B1(new_n810), .B2(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT89), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  OR2_X1    g391(.A1(G25), .A2(G29), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n816), .B2(new_n817), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n688), .A2(G24), .ZN(new_n822));
  INV_X1    g397(.A(G290), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n688), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1986), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n820), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n807), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n807), .A2(new_n826), .A3(KEYINPUT90), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(KEYINPUT34), .B1(new_n802), .B2(new_n806), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n793), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n793), .A3(new_n832), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n792), .B1(new_n834), .B2(new_n835), .ZN(G311));
  AND3_X1   g411(.A1(new_n791), .A2(new_n781), .A3(new_n708), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n831), .A2(new_n793), .A3(new_n832), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n837), .B(new_n706), .C1(new_n838), .C2(new_n833), .ZN(G150));
  NAND2_X1  g414(.A1(new_n606), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT101), .B(G93), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n522), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n545), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n525), .A2(G55), .B1(new_n846), .B2(G651), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n561), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n556), .A2(new_n560), .B1(new_n843), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n841), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n854), .B2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n848), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(G145));
  XOR2_X1   g435(.A(new_n487), .B(G160), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n631), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n773), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n502), .B(new_n755), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n773), .B(KEYINPUT103), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n723), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n866), .A2(new_n772), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n866), .A2(new_n772), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(new_n722), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(G130), .A2(new_n482), .B1(new_n466), .B2(G142), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n879), .A2(new_n481), .A3(G118), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n481), .B2(G118), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT105), .ZN(new_n884));
  INV_X1    g459(.A(new_n619), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n815), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n884), .A2(new_n885), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT106), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT106), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n877), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n872), .B(new_n876), .C1(new_n891), .C2(new_n892), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n863), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n889), .A2(new_n890), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n862), .B1(new_n877), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(G37), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n897), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n897), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(new_n614), .B(new_n852), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n605), .A2(new_n905), .A3(new_n784), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n534), .A2(G92), .A3(new_n535), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n600), .B1(new_n909), .B2(new_n603), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n910), .B2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(G299), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT41), .A4(new_n912), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n918), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n904), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G303), .B(new_n823), .ZN(new_n922));
  XOR2_X1   g497(.A(G288), .B(G305), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n913), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n904), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n925), .B1(new_n921), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n848), .A2(new_n594), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(G295));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n932), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(G286), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(G168), .B1(new_n552), .B2(new_n553), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n851), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n851), .B1(new_n938), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n927), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n852), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n851), .A2(new_n938), .A3(new_n939), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n915), .A2(new_n916), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n949), .A3(KEYINPUT111), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n946), .A2(new_n945), .B1(new_n915), .B2(new_n916), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n917), .A2(new_n919), .A3(new_n947), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n942), .A2(new_n913), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n924), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n958), .ZN(new_n961));
  INV_X1    g536(.A(new_n924), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n955), .B1(new_n963), .B2(new_n959), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI211_X1 g541(.A(KEYINPUT110), .B(new_n955), .C1(new_n963), .C2(new_n959), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n935), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND4_X1   g543(.A1(KEYINPUT43), .A2(new_n954), .A3(new_n956), .A4(new_n959), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n963), .B2(new_n959), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  NOR4_X1   g548(.A1(new_n472), .A2(new_n473), .A3(new_n973), .A4(new_n478), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n502), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n773), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT113), .Z(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n755), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n980), .B2(new_n772), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n887), .A2(new_n819), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n815), .A2(new_n818), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n979), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  NAND2_X1  g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n978), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n974), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  INV_X1    g572(.A(new_n977), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n997), .B(new_n998), .C1(new_n502), .C2(new_n975), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n976), .A2(new_n977), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n997), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT56), .B(G2072), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n572), .A2(KEYINPUT120), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n572), .A2(KEYINPUT120), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n574), .A3(new_n575), .A4(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1007), .A2(new_n1008), .B1(KEYINPUT57), .B2(new_n784), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n502), .A2(new_n1012), .A3(new_n975), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n974), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n787), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1004), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n473), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(G40), .A3(new_n477), .A4(new_n471), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n976), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1014), .A2(new_n711), .B1(new_n983), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(new_n605), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1004), .A2(new_n1015), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1009), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1017), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1016), .A2(KEYINPUT61), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT61), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1004), .A2(new_n1010), .A3(new_n1027), .A4(new_n1015), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n502), .A2(new_n975), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1019), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n976), .A2(KEYINPUT114), .A3(new_n977), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1002), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT58), .B(G1341), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1033), .A2(G1996), .B1(new_n1020), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n562), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1035), .B2(new_n562), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1029), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1040), .B(new_n910), .C1(new_n1021), .C2(KEYINPUT60), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1020), .A2(new_n983), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1011), .A2(new_n974), .A3(new_n1013), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT60), .B(new_n1042), .C1(new_n1043), .C2(G1348), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n605), .B1(new_n1044), .B2(KEYINPUT122), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1041), .A2(new_n1045), .B1(KEYINPUT122), .B2(new_n1044), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1021), .A2(KEYINPUT60), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1025), .B1(new_n1039), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT126), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1018), .A2(G40), .A3(new_n471), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n476), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(G2105), .B1(new_n476), .B2(new_n1054), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1052), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n472), .A2(new_n473), .A3(new_n973), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1057), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(KEYINPUT125), .A3(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(G2078), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n976), .B2(new_n977), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n995), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1051), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(KEYINPUT126), .A3(new_n995), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1031), .A2(new_n1002), .A3(new_n739), .A4(new_n1032), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n1063), .B1(new_n1073), .B2(new_n1014), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1071), .A2(new_n1074), .A3(G301), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT118), .B(new_n974), .C1(new_n1030), .C2(KEYINPUT45), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n502), .B2(new_n975), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n1019), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1030), .A2(new_n998), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(new_n1065), .ZN(new_n1082));
  AOI21_X1  g657(.A(G301), .B1(new_n1082), .B2(new_n1074), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1050), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G303), .A2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT115), .B(G1971), .Z(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1014), .A2(G2090), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(G8), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1019), .B2(new_n976), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G1976), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1093), .B(new_n1095), .C1(new_n1094), .C2(G288), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G305), .A2(G1981), .ZN(new_n1097));
  INV_X1    g672(.A(G1981), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT116), .B(G86), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n522), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1100), .B2(new_n585), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT49), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1097), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(new_n1093), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(new_n1094), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT52), .B1(new_n1092), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1096), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1014), .A2(KEYINPUT117), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1011), .A2(new_n1111), .A3(new_n974), .A4(new_n1013), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1110), .A2(new_n749), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1088), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1033), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1091), .B(new_n1108), .C1(new_n1116), .C2(new_n1087), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1081), .A2(new_n702), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1043), .A2(new_n731), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(G286), .A2(G8), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT123), .Z(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1081), .A2(new_n702), .B1(new_n731), .B2(new_n1043), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1127), .A2(new_n1109), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1119), .B(new_n1124), .C1(new_n1127), .C2(new_n1109), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1084), .A2(new_n1118), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1082), .A2(new_n1074), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n1132), .B2(G171), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1133), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1049), .A2(new_n1131), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1127), .A2(new_n1109), .A3(G286), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1117), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(G8), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1087), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n1091), .A3(new_n1108), .A4(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1097), .B1(new_n1105), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n1092), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(new_n1108), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1125), .B1(new_n1122), .B2(G8), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT62), .B(new_n1130), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n1083), .A3(new_n1118), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT62), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1149), .B(new_n1154), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n994), .B1(new_n1140), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n978), .B1(new_n772), .B2(new_n984), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n978), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT46), .B1(new_n978), .B2(G1996), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT47), .Z(new_n1166));
  NOR2_X1   g741(.A1(new_n978), .A2(new_n991), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT48), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n990), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n986), .A2(new_n987), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n755), .A2(G2067), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n978), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1161), .A2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g749(.A1(new_n966), .A2(new_n967), .ZN(new_n1176));
  OR2_X1    g750(.A1(G227), .A2(new_n461), .ZN(new_n1177));
  NOR3_X1   g751(.A1(G229), .A2(G401), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g752(.A(new_n895), .ZN(new_n1179));
  INV_X1    g753(.A(new_n723), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n868), .B2(new_n870), .ZN(new_n1181));
  OAI21_X1  g755(.A(new_n898), .B1(new_n1181), .B2(new_n875), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(new_n863), .ZN(new_n1183));
  OAI21_X1  g757(.A(new_n956), .B1(new_n1179), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n1178), .B1(new_n1184), .B2(new_n896), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n1176), .A2(new_n1185), .ZN(G308));
  OAI221_X1 g760(.A(new_n1178), .B1(new_n896), .B2(new_n1184), .C1(new_n966), .C2(new_n967), .ZN(G225));
endmodule


