//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  OR2_X1    g0000(.A1(KEYINPUT64), .A2(G50), .ZN(new_n201));
  NAND2_X1  g0001(.A1(KEYINPUT64), .A2(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(G58), .A2(G68), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n215), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  INV_X1    g0026(.A(KEYINPUT1), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n205), .A2(G50), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n230), .A2(new_n213), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n215), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT0), .Z(new_n235));
  NOR4_X1   g0035(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G169), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT76), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT13), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT74), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n231), .ZN(new_n260));
  NAND3_X1  g0060(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT69), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n262), .A2(new_n266), .A3(new_n263), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n218), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT67), .B(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G45), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n256), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n262), .A2(new_n266), .A3(new_n263), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n278));
  OAI21_X1  g0078(.A(G238), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(KEYINPUT74), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n260), .A2(new_n257), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n238), .A2(G1698), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n288), .C1(G226), .C2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G97), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n282), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n255), .B1(new_n281), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g0095(.A(KEYINPUT13), .B(new_n293), .C1(new_n276), .C2(new_n280), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n254), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n268), .A2(new_n256), .A3(new_n275), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT74), .B1(new_n279), .B2(new_n274), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n281), .A2(new_n255), .A3(new_n294), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G179), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT14), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n231), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n212), .A2(G20), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(G68), .A3(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n312), .B(KEYINPUT75), .Z(new_n313));
  NOR2_X1   g0113(.A1(G20), .A2(G33), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n284), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G77), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n309), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT11), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n307), .A2(new_n217), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(KEYINPUT11), .A3(new_n309), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(KEYINPUT14), .B(new_n254), .C1(new_n295), .C2(new_n296), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n305), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(G200), .B1(new_n295), .B2(new_n296), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n301), .A2(G190), .A3(new_n302), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n327), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n282), .ZN(new_n335));
  INV_X1    g0135(.A(G223), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT3), .A2(G33), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  OAI21_X1  g0138(.A(G1698), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n287), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G222), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n345), .A2(new_n346), .B1(new_n318), .B2(new_n287), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n335), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(G226), .B1(new_n277), .B2(new_n278), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n274), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n253), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT8), .B(G58), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  INV_X1    g0153(.A(new_n314), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n352), .A2(new_n317), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT71), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(new_n206), .B2(new_n213), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT8), .B(G58), .Z(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n316), .B1(G150), .B2(new_n314), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(KEYINPUT71), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n309), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n310), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n311), .A2(G50), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n362), .A2(new_n363), .B1(G50), .B2(new_n306), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n350), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT72), .B1(new_n351), .B2(new_n366), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT73), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n351), .A2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n370), .A4(new_n367), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n352), .B1(new_n212), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n310), .B1(new_n307), .B2(new_n352), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n285), .A2(new_n213), .A3(new_n286), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n213), .A4(new_n286), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(G68), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G58), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n217), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n393), .B2(new_n204), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n314), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n309), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n217), .B1(new_n385), .B2(new_n387), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n396), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(KEYINPUT16), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n382), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n264), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G232), .B1(new_n271), .B2(new_n273), .ZN(new_n407));
  AOI21_X1  g0207(.A(G1698), .B1(new_n285), .B2(new_n286), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G223), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n287), .A2(G226), .A3(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n335), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n253), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n407), .A2(new_n413), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(G179), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT18), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n407), .A2(new_n413), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n419), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT16), .B1(new_n391), .B2(new_n397), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n337), .A2(new_n338), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT7), .B1(new_n424), .B2(new_n213), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n425), .B2(new_n389), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n309), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n381), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n418), .B1(new_n422), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G200), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n407), .B2(new_n413), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G190), .B2(new_n415), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n405), .A2(new_n433), .A3(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n419), .A2(G169), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n369), .B2(new_n419), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n417), .A2(new_n430), .A3(new_n434), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT9), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n366), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n361), .A2(KEYINPUT9), .A3(new_n365), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT10), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n368), .A2(G190), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n350), .A2(G200), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(new_n442), .A3(new_n447), .A4(new_n443), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n218), .B1(new_n340), .B2(new_n342), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n424), .A2(G107), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n345), .B2(new_n238), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n335), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G244), .B1(new_n277), .B2(new_n278), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n274), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G200), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n307), .A2(new_n318), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n311), .A2(G77), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n362), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n358), .A2(new_n314), .B1(G20), .B2(G77), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT15), .B(G87), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n317), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n464), .B2(new_n309), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n455), .A2(G190), .A3(new_n274), .A4(new_n456), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n458), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n456), .A2(new_n274), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n340), .A2(new_n342), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G238), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n408), .A2(G232), .B1(new_n424), .B2(G107), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n282), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n253), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n455), .A2(new_n369), .A3(new_n274), .A4(new_n456), .ZN(new_n474));
  INV_X1    g0274(.A(new_n465), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n467), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n379), .A2(new_n440), .A3(new_n451), .A4(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n306), .A2(G116), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n212), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n306), .A2(new_n482), .A3(new_n231), .A4(new_n308), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n284), .B2(G97), .ZN(new_n486));
  NAND3_X1  g0286(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n308), .A2(new_n231), .B1(G20), .B2(new_n484), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n485), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G264), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n497));
  OAI211_X1 g0297(.A(G257), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n285), .A2(G303), .A3(new_n286), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n335), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n270), .A2(G1), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  OR2_X1    g0303(.A1(new_n503), .A2(G41), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n502), .B(new_n504), .C1(new_n269), .C2(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G270), .A3(new_n262), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n506), .A3(G179), .ZN(new_n507));
  XOR2_X1   g0307(.A(KEYINPUT67), .B(G41), .Z(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(G274), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n509), .A2(new_n262), .A3(new_n504), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n496), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n501), .A2(new_n506), .A3(new_n512), .ZN(new_n515));
  INV_X1    g0315(.A(new_n483), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n480), .B1(new_n516), .B2(G116), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n490), .A2(KEYINPUT20), .A3(new_n491), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n490), .B2(new_n491), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n520), .A3(G169), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT21), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n515), .A2(new_n520), .A3(new_n523), .A4(G169), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n514), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n335), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n505), .A2(G264), .A3(new_n262), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n512), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n253), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n213), .B2(G107), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT23), .A3(G20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n284), .A2(new_n484), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n213), .ZN(new_n540));
  AND2_X1   g0340(.A1(KEYINPUT83), .A2(G87), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n213), .B(new_n541), .C1(new_n337), .C2(new_n338), .ZN(new_n542));
  AND2_X1   g0342(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n543));
  NOR2_X1   g0343(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n538), .B(new_n540), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(new_n285), .B2(new_n286), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT24), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n547), .A3(new_n541), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n545), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n535), .A2(new_n537), .B1(new_n539), .B2(new_n213), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n401), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n536), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n306), .B2(G107), .ZN(new_n559));
  AOI22_X1  g0359(.A1(G107), .A2(new_n516), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  OAI221_X1 g0361(.A(new_n533), .B1(G179), .B2(new_n532), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n550), .A2(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n309), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n530), .A2(new_n531), .A3(new_n512), .A4(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n532), .A2(G200), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n564), .A2(new_n560), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n520), .B1(new_n515), .B2(G200), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n421), .B2(new_n515), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n525), .A2(new_n562), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n505), .A2(G257), .A3(new_n262), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n572), .A2(new_n512), .ZN(new_n573));
  INV_X1    g0373(.A(new_n489), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n487), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT4), .B1(new_n408), .B2(G244), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n335), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n573), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n581), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n572), .A2(new_n512), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT80), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n572), .A2(new_n512), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n582), .B1(new_n588), .B2(new_n369), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n306), .A2(G97), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n516), .B2(G97), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n388), .A2(G107), .A3(new_n390), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n290), .A2(new_n536), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G97), .A2(G107), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n536), .A2(KEYINPUT6), .A3(G97), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(G20), .B1(G77), .B2(new_n314), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT78), .B1(new_n600), .B2(new_n309), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT78), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n602), .B(new_n401), .C1(new_n592), .C2(new_n599), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n591), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n581), .A2(G190), .A3(new_n572), .A4(new_n512), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT81), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT81), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n573), .A2(new_n608), .A3(G190), .A4(new_n581), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(new_n309), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n602), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n309), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n572), .A2(new_n512), .A3(new_n586), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n586), .B1(new_n572), .B2(new_n512), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n581), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n610), .A2(new_n614), .A3(new_n591), .A4(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n213), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n219), .A2(new_n290), .A3(new_n536), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n213), .B(G68), .C1(new_n337), .C2(new_n338), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT19), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n623), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n309), .ZN(new_n629));
  INV_X1    g0429(.A(new_n463), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n306), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n516), .A2(KEYINPUT82), .A3(new_n630), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT82), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n483), .B2(new_n463), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n629), .A2(new_n632), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(G244), .B(G1698), .C1(new_n337), .C2(new_n338), .ZN(new_n637));
  OAI211_X1 g0437(.A(G238), .B(new_n344), .C1(new_n337), .C2(new_n338), .ZN(new_n638));
  INV_X1    g0438(.A(new_n539), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n335), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n510), .B1(new_n502), .B2(new_n220), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n262), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n369), .A3(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n640), .A2(new_n335), .B1(new_n642), .B2(new_n262), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n636), .B(new_n644), .C1(G169), .C2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n621), .A2(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n401), .B1(new_n647), .B2(new_n624), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n483), .A2(new_n219), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n631), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n641), .A2(G190), .A3(new_n643), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(new_n431), .C2(new_n645), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n571), .A2(new_n605), .A3(new_n619), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n334), .A2(new_n479), .A3(new_n654), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n430), .A2(new_n434), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n476), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n465), .B1(new_n457), .B2(new_n253), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(KEYINPUT85), .A3(new_n474), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n333), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n656), .B1(new_n330), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n417), .A2(new_n438), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n451), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n379), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n334), .A2(new_n479), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n589), .A2(new_n604), .A3(new_n653), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n589), .A2(new_n604), .A3(new_n653), .A4(KEYINPUT26), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n564), .A2(new_n560), .A3(new_n565), .A4(new_n566), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n525), .B2(new_n562), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(new_n619), .A3(new_n605), .A4(new_n653), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n676), .A3(new_n646), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n667), .A2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n212), .A2(new_n213), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n520), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n525), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n569), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n685), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n564), .B2(new_n560), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n562), .B1(new_n674), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n562), .A2(new_n685), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n525), .A2(new_n685), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n694), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n233), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n508), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n622), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n230), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT86), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n654), .B2(new_n685), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n618), .A2(new_n607), .A3(new_n609), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n605), .B(new_n653), .C1(new_n604), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n570), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT86), .A3(new_n691), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n583), .A2(new_n584), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n532), .A2(new_n507), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n645), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT30), .A4(new_n645), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n645), .A2(G179), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n617), .A2(new_n515), .A3(new_n532), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n685), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT31), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n710), .B1(new_n717), .B2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT87), .B(KEYINPUT29), .Z(new_n730));
  NAND3_X1  g0530(.A1(new_n677), .A2(new_n691), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n677), .A2(new_n691), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT87), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n729), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n709), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(G13), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n212), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n704), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n231), .B1(G20), .B2(new_n253), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n213), .A2(new_n369), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G190), .A3(new_n431), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n287), .B1(new_n747), .B2(new_n219), .C1(new_n392), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n421), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G50), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n755), .A2(KEYINPUT32), .A3(new_n756), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n213), .A2(new_n431), .A3(G179), .A4(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G107), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT32), .B1(new_n755), .B2(new_n756), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n753), .A2(new_n757), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n748), .A2(new_n754), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(KEYINPUT89), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n750), .B(new_n761), .C1(G77), .C2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n421), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n213), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n751), .A2(G190), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT90), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(KEYINPUT90), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n767), .B(new_n771), .C1(new_n217), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n775), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n749), .A2(new_n780), .B1(new_n762), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n755), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n287), .B(new_n782), .C1(G329), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n769), .ZN(new_n785));
  INV_X1    g0585(.A(new_n747), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G294), .B1(new_n786), .B2(G303), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n752), .A2(G326), .B1(G283), .B2(new_n758), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n779), .A2(new_n784), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n745), .B1(new_n776), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n745), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT88), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n251), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n703), .A2(new_n287), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G45), .C2(new_n230), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n233), .A2(new_n287), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n800), .B1(G116), .B2(new_n233), .C1(new_n210), .C2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n743), .B(new_n790), .C1(new_n797), .C2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n689), .B2(new_n794), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT92), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n688), .A2(new_n710), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n690), .A2(new_n743), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT93), .ZN(G396));
  AOI21_X1  g0609(.A(KEYINPUT86), .B1(new_n715), .B2(new_n691), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n714), .A2(new_n711), .A3(new_n570), .A4(new_n685), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n728), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G330), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n465), .A2(new_n691), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(new_n658), .B2(new_n660), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n814), .B1(new_n467), .B2(new_n476), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT96), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n659), .A2(KEYINPUT85), .A3(new_n474), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT85), .B1(new_n659), .B2(new_n474), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT96), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n477), .A2(new_n815), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n732), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n825), .A2(new_n677), .A3(new_n691), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n742), .B1(new_n813), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n813), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n744), .A2(new_n791), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n742), .B1(G77), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n749), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(G294), .B1(new_n783), .B2(G311), .ZN(new_n836));
  INV_X1    g0636(.A(new_n758), .ZN(new_n837));
  INV_X1    g0637(.A(G303), .ZN(new_n838));
  INV_X1    g0638(.A(new_n752), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n836), .B1(new_n219), .B2(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(G116), .B2(new_n766), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT94), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n287), .B1(new_n786), .B2(G107), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n777), .A2(G283), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(new_n842), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n844), .A3(new_n771), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n785), .A2(G58), .B1(new_n786), .B2(G50), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n424), .B1(new_n783), .B2(G132), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(new_n217), .C2(new_n837), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT95), .Z(new_n850));
  AOI22_X1  g0650(.A1(G137), .A2(new_n752), .B1(new_n835), .B2(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n851), .B1(new_n756), .B2(new_n765), .C1(new_n775), .C2(new_n353), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n846), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n834), .B1(new_n857), .B2(new_n744), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n825), .B2(new_n792), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n831), .A2(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n739), .A2(new_n212), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n327), .A2(new_n691), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT97), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n297), .A2(new_n303), .A3(new_n304), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n329), .A2(new_n328), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n333), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n330), .B2(new_n333), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n399), .B1(new_n402), .B2(new_n396), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n404), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n683), .B1(new_n871), .B2(new_n381), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n439), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n416), .A2(new_n683), .B1(new_n381), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n422), .A2(new_n429), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n405), .A2(new_n433), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n436), .A2(new_n429), .ZN(new_n878));
  INV_X1    g0678(.A(new_n683), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n429), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n877), .A2(new_n878), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n873), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n873), .A2(new_n883), .A3(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n869), .A2(new_n812), .A3(new_n825), .A4(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT40), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n826), .B1(new_n717), .B2(new_n728), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT98), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n439), .A2(new_n429), .A3(new_n879), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n882), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n439), .A2(new_n872), .B1(new_n876), .B2(new_n882), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT98), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n894), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n892), .A2(new_n903), .A3(KEYINPUT40), .A4(new_n869), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n891), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n812), .A2(new_n668), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n710), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n906), .B2(new_n905), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(KEYINPUT98), .A3(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n887), .A2(new_n893), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n910), .C1(new_n911), .C2(new_n899), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n886), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n330), .A2(new_n685), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n663), .A2(new_n683), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n659), .A2(new_n474), .A3(new_n691), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n828), .A2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n869), .A2(new_n920), .A3(new_n888), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n916), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n735), .A2(new_n668), .A3(new_n731), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT99), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT99), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n735), .A2(new_n668), .A3(new_n925), .A4(new_n731), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n666), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n922), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n861), .B1(new_n908), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n908), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n598), .A2(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n598), .A2(KEYINPUT35), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n231), .A2(new_n213), .A3(new_n484), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT36), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n230), .A2(new_n318), .A3(new_n393), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n203), .A2(new_n217), .ZN(new_n937));
  OAI211_X1 g0737(.A(G1), .B(new_n738), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n935), .A3(new_n938), .ZN(G367));
  NAND2_X1  g0739(.A1(new_n799), .A2(new_n244), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n795), .B1(new_n703), .B2(new_n630), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n743), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n650), .A2(new_n691), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n653), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n646), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n777), .A2(G294), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n769), .A2(new_n536), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n837), .A2(new_n290), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(G311), .C2(new_n752), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n424), .B1(new_n755), .B2(new_n951), .C1(new_n749), .C2(new_n838), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n747), .A2(new_n484), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(KEYINPUT46), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(KEYINPUT46), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n766), .B2(G283), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n947), .A2(new_n950), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n777), .A2(G159), .B1(new_n203), .B2(new_n766), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT103), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n770), .A2(G68), .ZN(new_n961));
  INV_X1    g0761(.A(G137), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n287), .B1(new_n755), .B2(new_n962), .C1(new_n749), .C2(new_n353), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n752), .A2(G143), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n318), .B2(new_n837), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n963), .B(new_n965), .C1(G58), .C2(new_n786), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n961), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n958), .A2(new_n959), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n957), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT47), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n942), .B1(new_n794), .B2(new_n946), .C1(new_n970), .C2(new_n745), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT101), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n605), .A2(new_n691), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n604), .A2(new_n685), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n619), .A2(new_n605), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT100), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT100), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n699), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT42), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n978), .A2(KEYINPUT101), .A3(KEYINPUT42), .A4(new_n699), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  INV_X1    g0784(.A(new_n946), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n976), .A2(new_n977), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n605), .B1(new_n986), .B2(new_n562), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n691), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n980), .B2(new_n979), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n985), .A2(new_n984), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n981), .A2(new_n982), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n989), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n697), .A2(new_n978), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT102), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(KEYINPUT102), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n991), .A2(new_n997), .A3(new_n995), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n704), .B(KEYINPUT41), .Z(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n973), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n986), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1008), .B2(new_n701), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n978), .A2(KEYINPUT44), .A3(new_n700), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(KEYINPUT45), .A3(new_n701), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n978), .B2(new_n700), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n696), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n695), .B(new_n698), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(new_n690), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1011), .A2(new_n697), .A3(new_n1015), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n736), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1005), .B1(new_n1021), .B2(new_n736), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1004), .B1(new_n1022), .B2(new_n741), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n971), .B1(new_n1003), .B2(new_n1023), .ZN(G387));
  INV_X1    g0824(.A(new_n762), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1025), .A2(G68), .B1(new_n783), .B2(G150), .ZN(new_n1026));
  INV_X1    g0826(.A(G50), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n287), .C1(new_n1027), .C2(new_n749), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n949), .B(new_n1028), .C1(G77), .C2(new_n786), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n752), .A2(G159), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT106), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n770), .A2(new_n630), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n777), .A2(new_n358), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n287), .B1(new_n783), .B2(G326), .ZN(new_n1035));
  INV_X1    g0835(.A(G283), .ZN(new_n1036));
  INV_X1    g0836(.A(G294), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n769), .A2(new_n1036), .B1(new_n747), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G322), .A2(new_n752), .B1(new_n835), .B2(G317), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n838), .B2(new_n765), .C1(new_n775), .C2(new_n781), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT49), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1035), .B1(new_n484), .B2(new_n837), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n744), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n801), .A2(new_n706), .B1(G107), .B2(new_n233), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n241), .A2(new_n270), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n706), .ZN(new_n1051));
  AOI211_X1 g0851(.A(G45), .B(new_n1051), .C1(G68), .C2(G77), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n352), .A2(G50), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n703), .B(new_n287), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1049), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT105), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n797), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1048), .B(new_n742), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n695), .B2(new_n793), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1019), .A2(new_n741), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT104), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(KEYINPUT104), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n736), .A2(new_n1019), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n704), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n736), .A2(new_n1019), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n978), .A2(new_n793), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT107), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n799), .A2(new_n248), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n795), .B1(G97), .B2(new_n703), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT108), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(KEYINPUT108), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n742), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n839), .A2(new_n951), .B1(new_n781), .B2(new_n749), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n759), .B1(new_n1036), .B2(new_n747), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n424), .B1(new_n755), .B2(new_n780), .C1(new_n1037), .C2(new_n762), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G116), .C2(new_n785), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(new_n838), .C2(new_n775), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT110), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n424), .B1(new_n783), .B2(G143), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n217), .B2(new_n747), .C1(new_n219), .C2(new_n837), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n358), .B2(new_n766), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n777), .A2(new_n203), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n770), .A2(G77), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G150), .A2(new_n752), .B1(new_n835), .B2(G159), .ZN(new_n1093));
  XOR2_X1   g0893(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1087), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1079), .B1(new_n1098), .B2(new_n744), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1073), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n740), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1067), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT111), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT111), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1105), .A3(new_n1067), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1021), .A2(new_n704), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  OAI21_X1  g0910(.A(new_n742), .B1(new_n358), .B2(new_n833), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n758), .A2(new_n203), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  INV_X1    g0913(.A(G132), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n287), .B1(new_n755), .B2(new_n1113), .C1(new_n749), .C2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(G128), .C2(new_n752), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n770), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1116), .B1(new_n962), .B2(new_n775), .C1(new_n756), .C2(new_n1117), .ZN(new_n1118));
  OR3_X1    g0918(.A1(new_n747), .A2(KEYINPUT53), .A3(new_n353), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT53), .B1(new_n747), .B2(new_n353), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1120), .C1(new_n765), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n777), .A2(G107), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n766), .A2(G97), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n747), .A2(new_n219), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n424), .B1(new_n749), .B2(new_n484), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G283), .C2(new_n752), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1123), .A2(new_n1092), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n837), .A2(new_n217), .B1(new_n755), .B2(new_n1037), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT113), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1118), .A2(new_n1122), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1111), .B1(new_n1131), .B2(new_n744), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n914), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n792), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT114), .Z(new_n1135));
  NAND4_X1  g0935(.A1(new_n869), .A2(new_n812), .A3(G330), .A4(new_n825), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n869), .A2(new_n920), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1137), .A2(new_n915), .A3(new_n903), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1137), .A2(new_n915), .B1(new_n913), .B2(new_n912), .ZN(new_n1139));
  OAI211_X1 g0939(.A(KEYINPUT112), .B(new_n1136), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n915), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n914), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(KEYINPUT112), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT112), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n892), .A2(new_n1144), .A3(G330), .A4(new_n869), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n915), .A3(new_n903), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1140), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1135), .B1(new_n741), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n812), .A2(G330), .A3(new_n825), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n828), .B(new_n919), .C1(new_n867), .C2(new_n868), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1150), .A2(new_n1137), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1137), .B2(new_n1151), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n924), .A2(new_n926), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n729), .A2(new_n668), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n667), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n927), .B(new_n1156), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1140), .A3(new_n1147), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n704), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1149), .A2(new_n1162), .ZN(G378));
  NAND3_X1  g0963(.A1(new_n891), .A2(G330), .A3(new_n904), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n451), .B1(new_n372), .B2(new_n371), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n366), .A2(new_n879), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1167), .B(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n891), .A2(new_n1169), .A3(new_n904), .A4(G330), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1171), .A2(new_n922), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n922), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1160), .B1(new_n1140), .B2(new_n1147), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1157), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n927), .A2(KEYINPUT117), .A3(new_n1156), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1177), .A2(KEYINPUT118), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT118), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1180), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT117), .B1(new_n927), .B2(new_n1156), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1183), .B1(new_n1159), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1176), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT118), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1159), .A2(new_n1183), .A3(new_n1186), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1175), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT120), .B1(new_n1194), .B2(KEYINPUT57), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1190), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1171), .A2(new_n922), .A3(new_n1172), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT119), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1175), .B2(new_n1198), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n705), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1191), .A2(new_n1195), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1170), .A2(new_n791), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n742), .B1(new_n203), .B2(new_n833), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n835), .A2(G128), .B1(new_n1025), .B2(G137), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1113), .B2(new_n839), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT116), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n747), .B2(new_n1121), .ZN(new_n1208));
  OR3_X1    g1008(.A1(new_n747), .A2(new_n1121), .A3(new_n1207), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n1114), .B2(new_n775), .C1(new_n353), .C2(new_n1117), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n758), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n837), .A2(new_n392), .B1(new_n318), .B2(new_n747), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n424), .B(new_n269), .C1(new_n755), .C2(new_n1036), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n749), .A2(new_n536), .B1(new_n762), .B2(new_n463), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n961), .B1(new_n484), .B2(new_n839), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT115), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1220), .B1(new_n290), .B2(new_n775), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1027), .B1(G33), .B2(G41), .C1(new_n508), .C2(new_n287), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1216), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1204), .B1(new_n1230), .B2(new_n744), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1176), .A2(new_n741), .B1(new_n1203), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1202), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT121), .ZN(G375));
  NAND2_X1  g1034(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1236), .A2(new_n1005), .A3(new_n1158), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1154), .A2(new_n740), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n791), .B1(new_n867), .B2(new_n868), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n833), .A2(G68), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n424), .B1(new_n755), .B2(new_n838), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n839), .A2(new_n1037), .B1(new_n747), .B2(new_n290), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G77), .C2(new_n758), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n536), .B2(new_n765), .C1(new_n484), .C2(new_n775), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1032), .B1(new_n1036), .B2(new_n749), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT122), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n839), .A2(new_n1114), .B1(new_n837), .B2(new_n392), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G159), .B2(new_n786), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n749), .A2(new_n962), .B1(new_n762), .B2(new_n353), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n424), .B(new_n1249), .C1(G128), .C2(new_n783), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n775), .A2(new_n1121), .B1(new_n1117), .B2(new_n1027), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n1244), .A2(new_n1246), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n745), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n743), .B(new_n1240), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1238), .B1(new_n1239), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(new_n1258), .ZN(G381));
  OAI211_X1 g1059(.A(new_n1109), .B(new_n971), .C1(new_n1023), .C2(new_n1003), .ZN(new_n1260));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G384), .A2(G378), .A3(G381), .A4(new_n1261), .ZN(new_n1262));
  OR3_X1    g1062(.A1(G375), .A2(new_n1260), .A3(new_n1262), .ZN(G407));
  NOR2_X1   g1063(.A1(G375), .A2(G378), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(new_n1265), .C2(G343), .ZN(G409));
  NAND3_X1  g1066(.A1(new_n1202), .A2(G378), .A3(new_n1232), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1200), .A2(new_n741), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1203), .A2(new_n1231), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1188), .A2(new_n1005), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1162), .B(new_n1149), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n684), .A2(G213), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1160), .A2(KEYINPUT60), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(new_n1236), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n705), .B1(new_n1276), .B2(new_n1236), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n831), .A2(KEYINPUT124), .A3(new_n859), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1258), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G384), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1274), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1288), .A2(G2897), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1287), .B(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1275), .B2(new_n1287), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G387), .A2(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1260), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1261), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1261), .B2(new_n1298), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1295), .A2(new_n1260), .A3(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1288), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1287), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1292), .A2(new_n1294), .A3(new_n1305), .A4(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1306), .A2(new_n1310), .A3(new_n1307), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1306), .B2(new_n1290), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1304), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1301), .B1(new_n1295), .B2(new_n1260), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT126), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1309), .B1(new_n1315), .B2(new_n1321), .ZN(G405));
  OAI21_X1  g1122(.A(new_n1307), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1318), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1303), .A2(KEYINPUT126), .A3(new_n1304), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1287), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1233), .A2(G378), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1265), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1328), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1323), .B(new_n1326), .C1(new_n1264), .C2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(G402));
endmodule


