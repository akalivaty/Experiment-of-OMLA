//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n453, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n590, new_n593, new_n595, new_n596, new_n597, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g029(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n472), .B2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n472), .A2(G136), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n471), .A2(new_n463), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n468), .A2(new_n470), .A3(G138), .A4(new_n463), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .A4(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(G126), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n491), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT71), .B1(new_n497), .B2(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT6), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n498), .A2(new_n501), .B1(new_n497), .B2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(G88), .A3(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n498), .A2(new_n501), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n497), .A2(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(G543), .A3(new_n512), .ZN(new_n513));
  OAI221_X1 g088(.A(new_n508), .B1(new_n509), .B2(new_n500), .C1(new_n510), .C2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n511), .A2(new_n512), .A3(new_n507), .ZN(new_n518));
  INV_X1    g093(.A(G89), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(new_n513), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n522), .A2(G51), .B1(G63), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  NAND2_X1  g101(.A1(new_n522), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(new_n518), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G90), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n500), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n513), .B1(new_n518), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n537), .A2(new_n538), .A3(new_n500), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n537), .B2(new_n500), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT74), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n513), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n502), .A2(new_n552), .A3(G53), .A4(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n502), .A2(G91), .A3(new_n507), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n505), .B2(new_n506), .ZN(new_n557));
  AND2_X1   g132(.A1(G78), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n554), .A2(new_n560), .ZN(G299));
  OAI21_X1  g136(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n528), .A2(G87), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n522), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  NAND3_X1  g141(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n511), .A2(G86), .A3(new_n512), .A4(new_n507), .ZN(new_n568));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n505), .B2(new_n506), .ZN(new_n570));
  AND2_X1   g145(.A1(G73), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(G305));
  NAND2_X1  g148(.A1(new_n522), .A2(G47), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n528), .A2(G85), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n500), .C2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  INV_X1    g153(.A(G54), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n579), .A2(new_n513), .B1(new_n580), .B2(new_n500), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n518), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n581), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n578), .B1(G868), .B2(new_n586), .ZN(G284));
  OAI21_X1  g162(.A(new_n578), .B1(G868), .B2(new_n586), .ZN(G321));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G299), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(G168), .B2(new_n589), .ZN(G297));
  OAI21_X1  g166(.A(new_n590), .B1(G168), .B2(new_n589), .ZN(G280));
  INV_X1    g167(.A(G559), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n586), .B1(new_n593), .B2(G860), .ZN(G148));
  NOR2_X1   g169(.A1(new_n541), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n586), .A2(new_n593), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(G868), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g173(.A(KEYINPUT78), .B(KEYINPUT11), .ZN(new_n599));
  XNOR2_X1  g174(.A(G323), .B(new_n599), .ZN(G282));
  NAND2_X1  g175(.A1(new_n472), .A2(G2104), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT13), .ZN(new_n603));
  INV_X1    g178(.A(G2100), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n472), .A2(G135), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n483), .A2(G123), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n463), .A2(G111), .ZN(new_n609));
  OAI21_X1  g184(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND3_X1  g187(.A1(new_n605), .A2(new_n606), .A3(new_n612), .ZN(G156));
  XNOR2_X1  g188(.A(G2427), .B(G2438), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n617), .A2(KEYINPUT14), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2451), .B(G2454), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2443), .B(G2446), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT79), .Z(new_n627));
  INV_X1    g202(.A(G14), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n624), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(G401));
  XNOR2_X1  g206(.A(G2067), .B(G2678), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT80), .ZN(new_n633));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2072), .B(G2078), .Z(new_n636));
  NOR3_X1   g211(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT18), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(KEYINPUT17), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n639), .A2(new_n634), .A3(new_n633), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n634), .B1(new_n633), .B2(new_n636), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(KEYINPUT81), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(KEYINPUT81), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n633), .B2(new_n639), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n638), .B(new_n640), .C1(new_n642), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XNOR2_X1  g222(.A(G1971), .B(G1976), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT20), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  NOR3_X1   g231(.A1(new_n650), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n650), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G229));
  NAND3_X1  g240(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT25), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n463), .ZN(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(G139), .C2(new_n472), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT92), .Z(new_n671));
  MUX2_X1   g246(.A(G33), .B(new_n671), .S(G29), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n442), .ZN(new_n673));
  MUX2_X1   g248(.A(G5), .B(G301), .S(G16), .Z(new_n674));
  INV_X1    g249(.A(G1961), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G32), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n472), .A2(G141), .ZN(new_n680));
  INV_X1    g255(.A(G105), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n464), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n483), .A2(G129), .ZN(new_n683));
  NAND3_X1  g258(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT26), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n679), .B1(new_n687), .B2(new_n678), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT93), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n678), .A2(G35), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G162), .B2(new_n678), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT29), .B(G2090), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT31), .B(G11), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT94), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(G28), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n678), .B1(new_n699), .B2(G28), .ZN(new_n701));
  OAI221_X1 g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .C1(new_n611), .C2(new_n678), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n678), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n472), .A2(G140), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n463), .A2(G116), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n483), .A2(G128), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n704), .B1(new_n713), .B2(new_n678), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n702), .B1(new_n714), .B2(G2067), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n689), .A2(new_n691), .ZN(new_n716));
  AND4_X1   g291(.A1(new_n692), .A2(new_n696), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n539), .A2(new_n540), .ZN(new_n718));
  INV_X1    g293(.A(new_n536), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT83), .B(G16), .Z(new_n721));
  MUX2_X1   g296(.A(new_n720), .B(G19), .S(new_n721), .Z(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1341), .Z(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(KEYINPUT24), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n678), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G160), .B2(new_n678), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2084), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n678), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n678), .ZN(new_n731));
  OAI22_X1  g306(.A1(new_n714), .A2(G2067), .B1(G2078), .B2(new_n731), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n729), .B(new_n732), .C1(G2078), .C2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(G21), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G286), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1966), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n717), .A2(new_n723), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n721), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT95), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  INV_X1    g318(.A(G4), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G16), .ZN(new_n745));
  INV_X1    g320(.A(new_n586), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G16), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(G1348), .Z(new_n748));
  NOR4_X1   g323(.A1(new_n677), .A2(new_n738), .A3(new_n743), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n678), .A2(G25), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n472), .A2(G131), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n483), .A2(G119), .ZN(new_n753));
  OR2_X1    g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n678), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT82), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G290), .B(G24), .S(new_n721), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1986), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G23), .B(G288), .S(G16), .Z(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT33), .B(G1976), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  MUX2_X1   g344(.A(G6), .B(G305), .S(G16), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT85), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT32), .B(G1981), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n767), .A2(new_n768), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n721), .A2(G22), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT88), .Z(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n721), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1971), .Z(new_n778));
  NAND4_X1  g353(.A1(new_n769), .A2(new_n773), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n780));
  OAI21_X1  g355(.A(new_n764), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n750), .B1(new_n788), .B2(new_n789), .ZN(G311));
  INV_X1    g365(.A(new_n789), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n783), .B2(new_n784), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n749), .B1(new_n791), .B2(new_n792), .ZN(G150));
  INV_X1    g368(.A(KEYINPUT98), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n720), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT99), .B1(new_n541), .B2(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n541), .A2(KEYINPUT98), .ZN(new_n799));
  INV_X1    g374(.A(G55), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n800), .A2(new_n513), .B1(new_n518), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n803), .A2(KEYINPUT97), .A3(new_n500), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT97), .B1(new_n803), .B2(new_n500), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n798), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n796), .A2(new_n797), .A3(new_n799), .A4(new_n806), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n586), .A2(G559), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n810), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n815));
  AOI21_X1  g390(.A(G860), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n806), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(KEYINPUT37), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(G145));
  XOR2_X1   g397(.A(G160), .B(new_n611), .Z(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G162), .Z(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n712), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n712), .A2(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n687), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n491), .A2(KEYINPUT101), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n488), .A2(new_n490), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n495), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n713), .A2(KEYINPUT102), .ZN(new_n835));
  INV_X1    g410(.A(new_n687), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n827), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n834), .B1(new_n830), .B2(new_n837), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n670), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n483), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n463), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n472), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(new_n602), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n757), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n830), .A2(new_n837), .ZN(new_n849));
  INV_X1    g424(.A(new_n495), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n488), .A2(new_n490), .A3(new_n832), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n832), .B1(new_n488), .B2(new_n490), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n671), .A3(new_n838), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n841), .A2(new_n848), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n848), .B1(new_n841), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n825), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT103), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(new_n825), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n856), .A2(new_n857), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n863), .B2(new_n824), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(KEYINPUT40), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT40), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(G395));
  OAI21_X1  g443(.A(KEYINPUT106), .B1(new_n806), .B2(G868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n810), .B(new_n596), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n586), .A2(G299), .A3(KEYINPUT104), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT104), .B1(new_n586), .B2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n586), .A2(G299), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n874), .B2(new_n870), .ZN(new_n880));
  XOR2_X1   g455(.A(G288), .B(G305), .Z(new_n881));
  XNOR2_X1  g456(.A(G166), .B(G290), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n589), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  MUX2_X1   g463(.A(KEYINPUT106), .B(new_n869), .S(new_n888), .Z(G295));
  MUX2_X1   g464(.A(KEYINPUT106), .B(new_n869), .S(new_n888), .Z(G331));
  INV_X1    g465(.A(new_n883), .ZN(new_n891));
  INV_X1    g466(.A(new_n874), .ZN(new_n892));
  XNOR2_X1  g467(.A(G286), .B(G301), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n810), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n809), .A3(new_n808), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n810), .A3(KEYINPUT107), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n877), .B1(new_n901), .B2(new_n876), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n874), .A2(KEYINPUT109), .A3(new_n875), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n902), .A2(new_n903), .B1(new_n895), .B2(new_n897), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n891), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n878), .A2(new_n876), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n907), .A3(new_n899), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n895), .A2(new_n874), .A3(new_n897), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n883), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n883), .B1(new_n908), .B2(new_n909), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g495(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n906), .C2(new_n912), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n915), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n912), .B2(new_n917), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n905), .A2(new_n919), .A3(new_n911), .A4(new_n910), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n926), .B(KEYINPUT43), .C1(new_n912), .C2(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n916), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n928), .ZN(G397));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n834), .B2(G1384), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n473), .A2(new_n477), .A3(G40), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(G290), .A2(G1986), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT48), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n933), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n937));
  INV_X1    g512(.A(new_n934), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n712), .A2(G2067), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n712), .A2(G2067), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n687), .B(G1996), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n757), .A2(new_n760), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n757), .A2(new_n760), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n935), .B(new_n939), .C1(new_n946), .C2(new_n933), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n936), .B1(new_n942), .B2(new_n687), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n933), .A2(KEYINPUT46), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT46), .B1(new_n933), .B2(new_n949), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n940), .B1(new_n954), .B2(new_n945), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n947), .B(new_n953), .C1(new_n933), .C2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n934), .A2(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n957), .B(new_n958), .Z(new_n959));
  OAI21_X1  g534(.A(new_n933), .B1(new_n959), .B2(new_n946), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n853), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n491), .B2(new_n495), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n932), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n966));
  AOI21_X1  g541(.A(G1348), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n932), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n853), .A2(new_n968), .A3(new_n963), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G2067), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT60), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n967), .B2(new_n970), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n586), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1956), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n962), .B1(new_n853), .B2(new_n963), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n968), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT57), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n980), .B(new_n981), .C1(new_n554), .C2(new_n560), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND2_X1  g558(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n984));
  AND4_X1   g559(.A1(new_n554), .A2(new_n560), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n853), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n932), .B1(new_n965), .B2(new_n930), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(new_n442), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n979), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n986), .B1(new_n979), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(KEYINPUT61), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n971), .A2(KEYINPUT60), .A3(new_n746), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n979), .A2(new_n991), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT61), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n986), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n975), .A2(new_n994), .A3(new_n995), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n949), .A3(new_n988), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT58), .B(G1341), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n969), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n541), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n720), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(KEYINPUT122), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT123), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1000), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n996), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n986), .B(KEYINPUT120), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n979), .A2(new_n1016), .A3(new_n991), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n586), .B1(new_n967), .B2(new_n970), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n992), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1015), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G286), .A2(G8), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n1025), .B2(KEYINPUT125), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n965), .A2(new_n930), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n931), .A2(new_n968), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n964), .A2(new_n966), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1027), .B(G8), .C1(new_n1035), .C2(G286), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1029), .A2(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1025), .B(new_n1026), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1035), .A2(new_n1040), .A3(G8), .A4(G286), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT124), .B1(new_n1037), .B2(new_n1025), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1036), .A2(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(G303), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G303), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2090), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n964), .A2(new_n1052), .A3(new_n966), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT112), .B(G1971), .Z(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n987), .B2(new_n988), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1051), .B(G8), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n563), .A2(G1976), .A3(new_n564), .A4(new_n565), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n969), .A2(new_n1058), .A3(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1062), .A2(G8), .A3(new_n969), .A4(new_n1058), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G305), .A2(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n567), .A2(new_n1065), .A3(new_n572), .A4(new_n568), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(G8), .B(new_n969), .C1(new_n1067), .C2(KEYINPUT49), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1064), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n1066), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1060), .B(new_n1063), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1057), .A2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n977), .A2(new_n978), .A3(G2090), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1076), .B2(new_n1055), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1051), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n931), .A2(new_n968), .A3(new_n987), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT126), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n853), .A2(new_n963), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n932), .B1(new_n1084), .B2(new_n930), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT126), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n987), .A4(new_n1081), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n987), .A2(new_n443), .A3(new_n988), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n964), .A2(new_n966), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1089), .A2(new_n1080), .B1(new_n1090), .B2(new_n675), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1085), .A2(new_n1028), .A3(new_n1081), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(G301), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT54), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1075), .B(new_n1079), .C1(new_n1092), .C2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1088), .A2(G301), .A3(new_n1091), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT54), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1043), .A2(new_n1096), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1075), .A2(new_n1079), .A3(new_n1097), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(KEYINPUT62), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1043), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1024), .A2(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1037), .A2(new_n1038), .A3(G286), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1075), .A2(new_n1079), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT63), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n969), .A2(G8), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1056), .A2(new_n1060), .A3(new_n1116), .A4(new_n1063), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n987), .A2(new_n988), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1054), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n964), .A2(new_n1052), .A3(new_n966), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1038), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT63), .B1(new_n1122), .B2(new_n1051), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1112), .A2(new_n1113), .B1(new_n1124), .B2(new_n1111), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1066), .B(KEYINPUT115), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G288), .A2(G1976), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1116), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1115), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1128), .A2(new_n1129), .B1(new_n1056), .B2(new_n1074), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1110), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1074), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(new_n1079), .A3(new_n1056), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1035), .A2(G8), .A3(G168), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1113), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1123), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1075), .A3(new_n1111), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(KEYINPUT116), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1131), .A2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT127), .B(new_n961), .C1(new_n1109), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1006), .A2(KEYINPUT122), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1012), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n999), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n992), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1021), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1105), .B(new_n1144), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1110), .B(new_n1130), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1154), .B(new_n1155), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1143), .B1(new_n1158), .B2(new_n960), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n956), .B1(new_n1142), .B2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g735(.A(new_n461), .ZN(new_n1162));
  NOR3_X1   g736(.A1(G229), .A2(new_n1162), .A3(G227), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1163), .A2(new_n630), .ZN(new_n1164));
  AOI21_X1  g738(.A(new_n1164), .B1(new_n862), .B2(new_n864), .ZN(new_n1165));
  AND3_X1   g739(.A1(new_n1165), .A2(new_n925), .A3(new_n927), .ZN(G308));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n925), .A3(new_n927), .ZN(G225));
endmodule


