//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT65), .A2(G146), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G143), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT0), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n188), .A2(G143), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT65), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT65), .A2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n201), .B2(G143), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(KEYINPUT0), .B2(G128), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT64), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n197), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n194), .A2(new_n197), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n210), .A2(new_n212), .A3(new_n216), .A4(new_n213), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n215), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT68), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n207), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n224), .A3(G116), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G119), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n225), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n225), .B2(new_n227), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n191), .A2(new_n236), .A3(G128), .A4(new_n193), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT66), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT66), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(new_n198), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n189), .A2(new_n190), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(new_n192), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n237), .B1(new_n241), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n213), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n209), .A2(G137), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n217), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n220), .A2(new_n235), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g066(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n220), .A2(new_n249), .ZN(new_n254));
  INV_X1    g068(.A(new_n235), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n251), .B1(new_n256), .B2(new_n250), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(KEYINPUT71), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT69), .A2(G953), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT69), .A2(G953), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G237), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(G210), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT29), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(G902), .B1(new_n259), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n235), .A4(new_n249), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n215), .A2(new_n217), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n207), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n249), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n255), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n252), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n268), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n220), .A2(KEYINPUT30), .A3(new_n249), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n274), .A2(new_n249), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n255), .C1(new_n280), .C2(KEYINPUT30), .ZN(new_n281));
  INV_X1    g095(.A(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n250), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n271), .B1(new_n284), .B2(KEYINPUT29), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G472), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n281), .A2(new_n250), .A3(new_n268), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n281), .A2(KEYINPUT31), .A3(new_n250), .A4(new_n268), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n282), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT70), .B1(new_n277), .B2(new_n282), .ZN(new_n295));
  OAI22_X1  g109(.A1(new_n290), .A2(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n277), .A2(new_n282), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n288), .A2(new_n289), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n301), .A2(new_n293), .B1(new_n302), .B2(new_n291), .ZN(new_n303));
  INV_X1    g117(.A(new_n297), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n286), .B1(new_n298), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT22), .B(G137), .Z(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT76), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n201), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n321));
  OR3_X1    g135(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G110), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT67), .B(G119), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G128), .ZN(new_n328));
  AOI22_X1  g142(.A1(G119), .A2(new_n240), .B1(new_n327), .B2(G128), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n325), .B(new_n328), .C1(new_n329), .C2(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n240), .A2(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT24), .B(G110), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n339));
  INV_X1    g153(.A(new_n328), .ZN(new_n340));
  OAI21_X1  g154(.A(G110), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n323), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT73), .A4(G146), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n321), .A2(new_n322), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n188), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n334), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n329), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n336), .B2(KEYINPUT74), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n313), .B1(new_n338), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n330), .A2(new_n335), .ZN(new_n353));
  INV_X1    g167(.A(new_n324), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(KEYINPUT75), .A3(new_n337), .A4(new_n350), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n312), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n351), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n311), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n307), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI221_X1 g178(.A(new_n307), .B1(KEYINPUT77), .B2(KEYINPUT25), .C1(new_n359), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT72), .B(G217), .ZN(new_n368));
  INV_X1    g182(.A(G234), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n359), .A2(new_n361), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(G902), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n367), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G214), .B1(G237), .B2(G902), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n375), .B(KEYINPUT81), .Z(new_n376));
  NAND2_X1  g190(.A1(new_n245), .A2(new_n316), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n202), .A2(new_n206), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n191), .A2(new_n197), .A3(new_n193), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(G125), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G224), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G953), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT7), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n377), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n377), .B2(new_n380), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(KEYINPUT79), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n394), .A2(G107), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n393), .A3(new_n395), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT80), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G101), .C1(KEYINPUT80), .C2(new_n391), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n225), .A2(new_n227), .A3(new_n232), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n222), .A2(new_n224), .A3(new_n406), .A4(G116), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G113), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT82), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n225), .A2(KEYINPUT5), .A3(new_n227), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n407), .A2(new_n411), .A3(G113), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n225), .A2(KEYINPUT5), .A3(new_n227), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n403), .B1(new_n414), .B2(new_n408), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(new_n402), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n405), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT8), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n385), .A2(new_n386), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT83), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n410), .A2(G113), .A3(new_n407), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n423), .A2(new_n403), .A3(new_n400), .A4(new_n402), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n397), .B1(new_n398), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n395), .B1(new_n388), .B2(new_n391), .ZN(new_n427));
  OAI21_X1  g241(.A(G101), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n430), .B(G101), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n234), .B2(new_n233), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n424), .B(new_n418), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n236), .B1(new_n201), .B2(G143), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n202), .B1(new_n434), .B2(new_n240), .ZN(new_n435));
  AOI21_X1  g249(.A(G125), .B1(new_n435), .B2(new_n237), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n378), .A2(G125), .A3(new_n379), .ZN(new_n437));
  OAI22_X1  g251(.A1(new_n436), .A2(new_n437), .B1(new_n383), .B2(new_n382), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n377), .A2(new_n380), .A3(new_n384), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n415), .A2(new_n416), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n411), .B1(new_n407), .B2(G113), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n414), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n404), .B1(new_n444), .B2(new_n412), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n419), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n441), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n422), .A2(new_n433), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n424), .B1(new_n429), .B2(new_n432), .ZN(new_n449));
  INV_X1    g263(.A(new_n418), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n433), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n453), .A3(new_n450), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n436), .A2(new_n437), .A3(new_n382), .ZN(new_n455));
  INV_X1    g269(.A(new_n382), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n456), .B1(new_n377), .B2(new_n380), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G210), .B1(G237), .B2(G902), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n448), .A2(new_n307), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n448), .A2(new_n462), .A3(new_n307), .A4(new_n459), .ZN(new_n463));
  INV_X1    g277(.A(new_n460), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT84), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(KEYINPUT85), .A2(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n459), .A2(new_n307), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(new_n462), .A3(new_n448), .A4(new_n465), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n376), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n192), .A2(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n476), .A2(new_n263), .A3(G214), .A4(new_n264), .ZN(new_n477));
  OR2_X1    g291(.A1(KEYINPUT69), .A2(G953), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n478), .A2(G214), .A3(new_n264), .A4(new_n260), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT18), .A2(G131), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n477), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n320), .B1(new_n188), .B2(new_n319), .ZN(new_n483));
  INV_X1    g297(.A(new_n480), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT87), .B1(new_n192), .B2(KEYINPUT86), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n472), .A2(G143), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n479), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n482), .B(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT89), .B(G104), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT90), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n477), .A2(new_n216), .A3(new_n480), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n489), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT17), .B(G131), .C1(new_n484), .C2(new_n488), .ZN(new_n499));
  AOI21_X1  g313(.A(G146), .B1(new_n321), .B2(new_n322), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n342), .B2(new_n323), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n344), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n491), .B(new_n495), .C1(new_n498), .C2(new_n502), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n490), .B(new_n216), .C1(new_n477), .C2(new_n480), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n482), .A2(new_n483), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n318), .B1(KEYINPUT88), .B2(KEYINPUT19), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n508));
  NOR2_X1   g322(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n315), .B(new_n317), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n201), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n323), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n489), .B2(new_n497), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n494), .B1(new_n506), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G475), .A2(G902), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n471), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  AOI211_X1 g332(.A(KEYINPUT20), .B(new_n518), .C1(new_n503), .C2(new_n514), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n491), .B1(new_n498), .B2(new_n502), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n494), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n521), .B2(new_n503), .ZN(new_n522));
  INV_X1    g336(.A(G475), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n517), .A2(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n240), .A2(G143), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT13), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n196), .A2(G143), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(G134), .B1(new_n529), .B2(new_n525), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n238), .A2(new_n239), .A3(new_n192), .ZN(new_n531));
  NOR4_X1   g345(.A1(new_n531), .A2(new_n526), .A3(new_n209), .A4(new_n528), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT91), .B1(new_n226), .B2(G122), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n534));
  INV_X1    g348(.A(G122), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(G116), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n533), .A2(new_n536), .B1(new_n226), .B2(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT92), .B(G107), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n530), .A2(new_n532), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n536), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n390), .B1(new_n542), .B2(KEYINPUT14), .ZN(new_n543));
  INV_X1    g357(.A(new_n537), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI221_X1 g359(.A(new_n542), .B1(KEYINPUT14), .B2(new_n390), .C1(G116), .C2(new_n535), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n209), .B1(new_n531), .B2(new_n528), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n525), .A2(G134), .A3(new_n529), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT9), .B(G234), .Z(new_n551));
  INV_X1    g365(.A(G953), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n551), .A2(new_n552), .A3(new_n368), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n541), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n307), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G478), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(KEYINPUT15), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n557), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(G952), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(G234), .B2(G237), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n307), .B(new_n263), .C1(G234), .C2(G237), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n524), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n551), .ZN(new_n567));
  OAI21_X1  g381(.A(G221), .B1(new_n567), .B2(G902), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT78), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n263), .A2(G227), .ZN(new_n571));
  XOR2_X1   g385(.A(G110), .B(G140), .Z(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n416), .A2(new_n435), .A3(new_n237), .ZN(new_n574));
  INV_X1    g388(.A(new_n237), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n196), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n191), .B2(new_n193), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n400), .B(new_n402), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n218), .A2(new_n219), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n215), .B2(new_n217), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n581), .A2(new_n582), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n245), .A2(KEYINPUT10), .A3(new_n400), .A4(new_n402), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n428), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n207), .A3(new_n431), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n218), .A2(new_n219), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n573), .B1(new_n584), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n586), .A2(new_n589), .A3(new_n587), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n580), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n573), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n593), .B(G469), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G469), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n584), .A2(new_n598), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n595), .B2(new_n591), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n600), .B(new_n307), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n600), .A2(new_n307), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n566), .A2(new_n570), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n306), .A2(new_n374), .A3(new_n470), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NOR2_X1   g423(.A1(new_n303), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n610), .A2(new_n611), .B1(new_n304), .B2(new_n303), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n570), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n433), .B1(new_n421), .B2(KEYINPUT83), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n441), .B1(new_n440), .B2(new_n446), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n307), .B(new_n459), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n464), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n461), .ZN(new_n619));
  INV_X1    g433(.A(new_n376), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n554), .A2(new_n622), .A3(new_n556), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n558), .A2(G902), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT93), .B1(new_n553), .B2(KEYINPUT94), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n541), .B2(new_n549), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n541), .A2(new_n627), .A3(new_n549), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT94), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n626), .B1(new_n629), .B2(new_n555), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n623), .B(new_n624), .C1(new_n630), .C2(new_n622), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT95), .B(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n557), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n524), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n621), .A2(new_n565), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n614), .A2(new_n374), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND2_X1  g454(.A1(new_n515), .A2(new_n516), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT20), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n515), .A2(new_n471), .A3(new_n516), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n521), .A2(new_n503), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n307), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(G475), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n565), .B(KEYINPUT97), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n647), .A3(new_n560), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n376), .B1(new_n618), .B2(new_n461), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n642), .A2(new_n643), .B1(new_n646), .B2(G475), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n560), .A4(new_n648), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n650), .A2(new_n654), .A3(KEYINPUT99), .A4(new_n651), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n374), .A3(new_n614), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NAND2_X1  g476(.A1(new_n367), .A2(new_n371), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n352), .A2(new_n358), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n311), .A2(KEYINPUT36), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NOR4_X1   g481(.A1(new_n666), .A2(new_n667), .A3(G902), .A4(new_n371), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n611), .B1(new_n296), .B2(new_n307), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n303), .A2(new_n304), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n668), .B1(new_n367), .B2(new_n371), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT100), .B1(new_n676), .B2(new_n612), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n607), .A2(new_n470), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(new_n562), .ZN(new_n682));
  INV_X1    g496(.A(new_n563), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(G900), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT101), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n652), .A2(new_n560), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT102), .B1(new_n621), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n560), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n524), .A3(new_n685), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n651), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT32), .B1(new_n303), .B2(new_n304), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n296), .A2(new_n287), .A3(new_n297), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n613), .B1(new_n696), .B2(new_n286), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n693), .A2(new_n697), .A3(new_n670), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  INV_X1    g513(.A(new_n613), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n685), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n652), .A2(new_n689), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n704), .A2(new_n620), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n281), .A2(new_n250), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n268), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n256), .A2(new_n250), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n307), .B1(new_n711), .B2(new_n268), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n696), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n463), .A2(new_n466), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(new_n469), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n467), .A2(new_n469), .A3(new_n719), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n707), .A2(new_n670), .A3(new_n715), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n192), .ZN(G45));
  NAND3_X1  g539(.A1(new_n634), .A2(new_n524), .A3(new_n686), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT105), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n634), .A2(new_n524), .A3(new_n728), .A4(new_n686), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n727), .A2(new_n651), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n697), .A2(new_n670), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  OAI21_X1  g546(.A(new_n307), .B1(new_n601), .B2(new_n602), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G469), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n570), .A3(new_n603), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(KEYINPUT106), .A3(new_n570), .A4(new_n603), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n306), .A2(new_n636), .A3(new_n739), .A4(new_n374), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND2_X1  g556(.A1(new_n372), .A2(new_n373), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n663), .A2(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n694), .A2(new_n695), .B1(G472), .B2(new_n285), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n659), .A2(new_n746), .A3(new_n739), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR2_X1   g562(.A1(new_n621), .A2(new_n735), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n670), .A2(new_n306), .A3(new_n566), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  AND3_X1   g565(.A1(new_n737), .A2(new_n648), .A3(new_n738), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n296), .A2(new_n307), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT107), .B(G472), .ZN(new_n754));
  OAI22_X1  g568(.A1(new_n290), .A2(new_n292), .B1(new_n259), .B2(new_n268), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n753), .A2(new_n754), .B1(new_n297), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n651), .A2(new_n706), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n752), .A2(new_n374), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  AND2_X1   g574(.A1(new_n727), .A2(new_n729), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n670), .A2(new_n761), .A3(new_n749), .A4(new_n756), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT108), .B(G125), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G27));
  NAND4_X1  g578(.A1(new_n716), .A2(new_n717), .A3(new_n469), .A4(new_n620), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n467), .A2(KEYINPUT109), .A3(new_n620), .A4(new_n469), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n700), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT110), .A4(new_n700), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n746), .A3(new_n761), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(KEYINPUT42), .A3(new_n746), .A4(new_n761), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n746), .A3(new_n690), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n581), .A2(new_n582), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n579), .A2(new_n583), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n597), .B1(new_n785), .B2(new_n591), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n596), .A2(new_n598), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n593), .B(KEYINPUT45), .C1(new_n596), .C2(new_n598), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n789), .A3(G469), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n605), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n603), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(KEYINPUT111), .ZN(new_n793));
  INV_X1    g607(.A(new_n790), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n604), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT111), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n791), .B2(new_n603), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n793), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n569), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(new_n701), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n767), .A2(new_n768), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n631), .A2(new_n633), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT43), .B1(new_n804), .B2(new_n524), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n652), .A2(new_n806), .A3(new_n634), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n612), .A2(new_n670), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n803), .B1(new_n808), .B2(KEYINPUT44), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n801), .B(new_n809), .C1(KEYINPUT44), .C2(new_n808), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n799), .B2(new_n569), .ZN(new_n814));
  INV_X1    g628(.A(new_n798), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(KEYINPUT46), .B2(new_n795), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n570), .B(new_n812), .C1(new_n816), .C2(new_n793), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n744), .A2(new_n761), .A3(new_n745), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n802), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND4_X1  g635(.A1(new_n652), .A2(new_n620), .A3(new_n634), .A4(new_n570), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n734), .A2(new_n603), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT113), .Z(new_n825));
  AOI211_X1 g639(.A(new_n822), .B(new_n825), .C1(KEYINPUT49), .C2(new_n823), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n374), .A3(new_n723), .A4(new_n715), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n757), .A2(new_n613), .A3(new_n685), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n676), .A3(new_n714), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n698), .A2(new_n731), .A3(new_n829), .A4(new_n762), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT115), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n670), .B(new_n697), .C1(new_n693), .C2(new_n730), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n762), .A4(new_n829), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n306), .A2(new_n374), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n836), .B(new_n687), .C1(new_n771), .C2(new_n772), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n755), .A2(new_n297), .ZN(new_n838));
  INV_X1    g652(.A(new_n754), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n610), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n676), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n761), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n771), .B2(new_n772), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n524), .A2(new_n560), .A3(new_n685), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n767), .A2(new_n768), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n745), .A2(new_n676), .A3(new_n613), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n767), .A2(new_n768), .A3(KEYINPUT114), .A4(new_n844), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n837), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n652), .A2(new_n560), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n635), .ZN(new_n853));
  INV_X1    g667(.A(new_n648), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n614), .A2(new_n374), .A3(new_n855), .A4(new_n470), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n679), .A2(new_n608), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n659), .A2(new_n746), .A3(new_n739), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n740), .A2(new_n759), .A3(new_n750), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n778), .A2(new_n835), .A3(new_n851), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(new_n831), .B2(new_n834), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT53), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n679), .A2(new_n608), .A3(new_n856), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n744), .A2(new_n840), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n737), .A2(new_n648), .A3(new_n738), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n757), .ZN(new_n869));
  INV_X1    g683(.A(new_n735), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n651), .A3(new_n566), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n745), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n867), .A2(new_n869), .B1(new_n872), .B2(new_n670), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n866), .A2(new_n740), .A3(new_n747), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n843), .ZN(new_n875));
  INV_X1    g689(.A(new_n850), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n780), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n865), .A2(new_n878), .A3(new_n879), .A4(new_n778), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n863), .A2(new_n880), .A3(KEYINPUT54), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n879), .B1(new_n861), .B2(new_n862), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT116), .B1(new_n858), .B2(new_n859), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n873), .A2(new_n885), .A3(new_n740), .A4(new_n747), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT53), .A2(new_n884), .A3(new_n866), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n865), .A2(new_n887), .A3(new_n778), .A4(new_n851), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n882), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n734), .A2(new_n569), .A3(new_n603), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n814), .A2(new_n817), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n805), .A2(new_n562), .A3(new_n807), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(new_n374), .A3(new_n756), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n803), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n696), .A2(new_n374), .A3(new_n562), .A4(new_n713), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n634), .A2(new_n524), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n870), .A3(new_n802), .A4(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n870), .A2(new_n892), .A3(new_n767), .A4(new_n768), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n841), .ZN(new_n900));
  XNOR2_X1  g714(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n735), .A2(new_n620), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n723), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n893), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n902), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n722), .B2(new_n721), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(KEYINPUT50), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n867), .A2(new_n906), .A3(new_n892), .A4(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n898), .A2(new_n900), .A3(new_n904), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n867), .A2(new_n906), .A3(new_n892), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n912), .A2(new_n901), .B1(new_n899), .B2(new_n841), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n909), .A4(new_n898), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n895), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n814), .A2(new_n817), .A3(new_n920), .A4(new_n890), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n921), .A3(new_n894), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n910), .A2(new_n917), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  INV_X1    g739(.A(new_n896), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n802), .A2(new_n870), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n635), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n867), .A2(new_n749), .A3(new_n892), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(G952), .A3(new_n552), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n925), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n899), .A2(new_n746), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT48), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n928), .A2(new_n930), .A3(new_n925), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n918), .A2(new_n924), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n881), .A2(new_n889), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n881), .A2(new_n889), .A3(new_n937), .A4(KEYINPUT121), .ZN(new_n941));
  OR2_X1    g755(.A1(G952), .A2(G953), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n827), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n827), .C1(new_n940), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G75));
  NOR2_X1   g762(.A1(new_n263), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n307), .B1(new_n882), .B2(new_n888), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G210), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n452), .A2(new_n454), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n458), .ZN(new_n955));
  XOR2_X1   g769(.A(KEYINPUT123), .B(KEYINPUT55), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT56), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n950), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT56), .B1(new_n952), .B2(KEYINPUT124), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(KEYINPUT124), .B2(new_n952), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(new_n957), .ZN(G51));
  NAND2_X1  g776(.A1(new_n882), .A2(new_n888), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT54), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n889), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n604), .B(KEYINPUT57), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n602), .B2(new_n601), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n951), .A2(new_n794), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n949), .B1(new_n968), .B2(new_n969), .ZN(G54));
  AND3_X1   g784(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n950), .B1(new_n971), .B2(new_n515), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n515), .B2(new_n971), .ZN(G60));
  INV_X1    g787(.A(new_n623), .ZN(new_n974));
  INV_X1    g788(.A(new_n630), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(KEYINPUT33), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n965), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n881), .A2(new_n889), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n976), .B1(new_n981), .B2(new_n979), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n980), .A2(new_n949), .A3(new_n982), .ZN(G63));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n882), .B2(new_n888), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n666), .A2(new_n667), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n950), .C1(new_n372), .C2(new_n986), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n564), .B2(new_n381), .ZN(new_n991));
  INV_X1    g805(.A(new_n263), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n860), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(G898), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n954), .B1(new_n994), .B2(new_n992), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n993), .B(new_n995), .Z(G69));
  AND2_X1   g810(.A1(new_n810), .A2(new_n820), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n832), .A2(new_n762), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n836), .A2(new_n757), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n837), .B(new_n998), .C1(new_n801), .C2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n997), .A2(new_n778), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n263), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n279), .B1(new_n280), .B2(KEYINPUT30), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n507), .A2(new_n510), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(G900), .B2(new_n992), .ZN(new_n1006));
  OR4_X1    g820(.A1(new_n836), .A2(new_n803), .A3(new_n702), .A4(new_n853), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n724), .A2(KEYINPUT62), .A3(new_n998), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT62), .B1(new_n724), .B2(new_n998), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n997), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n263), .ZN(new_n1011));
  AOI22_X1  g825(.A1(new_n1002), .A2(new_n1006), .B1(new_n1011), .B2(new_n1005), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1012), .A2(KEYINPUT127), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1011), .A2(new_n1005), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1019), .B2(new_n1013), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1012), .A2(KEYINPUT126), .A3(new_n1014), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT126), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1022));
  OAI22_X1  g836(.A1(new_n1015), .A2(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(G72));
  NAND2_X1  g837(.A1(new_n1001), .A2(new_n860), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  AOI21_X1  g840(.A(new_n283), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1026), .B1(new_n1010), .B2(new_n874), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n710), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n950), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n863), .A2(new_n880), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n709), .A2(new_n283), .A3(new_n1026), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n1027), .B(new_n1030), .C1(new_n1031), .C2(new_n1032), .ZN(G57));
endmodule


