//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n201), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(KEYINPUT67), .A2(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(KEYINPUT67), .A2(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT68), .ZN(new_n233));
  INV_X1    g0033(.A(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  AND3_X1   g0036(.A1(new_n220), .A2(new_n235), .A3(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XOR2_X1   g0044(.A(G264), .B(G270), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(G222), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(G1698), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n261), .B1(new_n203), .B2(new_n259), .C1(new_n262), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n270), .A2(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n274), .A2(G226), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n268), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT72), .B(G200), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n284), .B2(new_n280), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n214), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT70), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n214), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n271), .A2(G13), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n215), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n271), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G50), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n215), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(G150), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n215), .A2(new_n256), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n215), .B1(new_n201), .B2(new_n202), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G13), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n296), .B(new_n303), .C1(G50), .C2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n285), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n285), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n280), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n307), .B1(new_n314), .B2(G169), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n280), .A2(G179), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G58), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT8), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT8), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n295), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n294), .A2(new_n325), .B1(new_n293), .B2(new_n297), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT66), .A2(G68), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT66), .A2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(G58), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n221), .A2(new_n332), .A3(G58), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n333), .A3(new_n217), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  INV_X1    g0135(.A(new_n300), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G159), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n257), .A2(new_n215), .A3(new_n258), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n258), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n221), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n337), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n287), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n334), .A2(G20), .B1(G159), .B2(new_n336), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n342), .B2(G68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n327), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(G223), .A2(G1698), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n352), .B1(G226), .B2(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n270), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n278), .A2(new_n270), .A3(G274), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n239), .B2(new_n273), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G179), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(new_n358), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT18), .B1(new_n351), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n349), .A2(new_n335), .A3(new_n337), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n287), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT16), .B1(new_n348), .B2(new_n343), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n326), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n361), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n355), .A2(new_n357), .A3(new_n281), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n355), .A2(new_n357), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(G200), .B2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n326), .C1(new_n365), .C2(new_n366), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n351), .A2(KEYINPUT17), .A3(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  OR3_X1    g0179(.A1(new_n306), .A2(KEYINPUT12), .A3(G68), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT12), .B1(new_n306), .B2(new_n221), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n381), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n298), .ZN(new_n386));
  AOI22_X1  g0186(.A1(G50), .A2(new_n336), .B1(new_n386), .B2(G77), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n215), .B2(new_n221), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n291), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n388), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n293), .A2(new_n287), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(G68), .A3(new_n295), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n385), .A2(new_n391), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G226), .A2(G1698), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n239), .B2(G1698), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n259), .B1(G33), .B2(G97), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n270), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n239), .A2(G1698), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G226), .B2(G1698), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n263), .A2(new_n264), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G238), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n356), .B1(new_n410), .B2(new_n273), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n397), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g0213(.A(KEYINPUT13), .B(new_n411), .C1(new_n402), .C2(new_n408), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n396), .B(G169), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n408), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT74), .B1(new_n407), .B2(new_n267), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(new_n397), .A3(new_n412), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(G179), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n420), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n396), .B1(new_n423), .B2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n395), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n395), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n413), .B2(new_n414), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(G190), .A3(new_n420), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(G232), .B(new_n260), .C1(new_n263), .C2(new_n264), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n257), .A2(G107), .A3(new_n258), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n265), .C2(new_n225), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n267), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n274), .A2(G244), .B1(new_n275), .B2(new_n278), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n360), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n215), .A2(new_n203), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(KEYINPUT71), .C1(new_n297), .C2(new_n300), .ZN(new_n440));
  XOR2_X1   g0240(.A(KEYINPUT15), .B(G87), .Z(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n386), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n323), .A2(new_n336), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT71), .B1(new_n444), .B2(new_n439), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n287), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n347), .A2(new_n306), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n295), .A2(G77), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n447), .A2(new_n448), .B1(G77), .B2(new_n306), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n437), .A2(new_n451), .A3(KEYINPUT73), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT73), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT71), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n300), .B1(new_n320), .B2(new_n322), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n438), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n442), .A3(new_n440), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n449), .B1(new_n457), .B2(new_n287), .ZN(new_n458));
  AOI21_X1  g0258(.A(G169), .B1(new_n434), .B2(new_n435), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n434), .A2(new_n435), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n436), .A2(new_n284), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n458), .C1(new_n281), .C2(new_n436), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NOR4_X1   g0266(.A1(new_n318), .A2(new_n379), .A3(new_n430), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT7), .B1(new_n406), .B2(new_n215), .ZN(new_n469));
  INV_X1    g0269(.A(new_n341), .ZN(new_n470));
  OAI21_X1  g0270(.A(G107), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n300), .A2(new_n203), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT6), .ZN(new_n473));
  AND2_X1   g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n206), .ZN(new_n475));
  INV_X1    g0275(.A(G107), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n472), .B1(new_n478), .B2(G20), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n347), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n306), .A2(G97), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n271), .A2(G33), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n289), .A2(new_n290), .A3(new_n306), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n480), .A2(KEYINPUT77), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT77), .ZN(new_n488));
  INV_X1    g0288(.A(new_n472), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n476), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n473), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(new_n215), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n476), .B1(new_n340), .B2(new_n341), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n287), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND4_X1   g0295(.A1(new_n289), .A2(new_n290), .A3(new_n306), .A4(new_n483), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n481), .B1(new_n496), .B2(G97), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n488), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n487), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G244), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G1698), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(new_n263), .B2(new_n264), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT78), .B1(G33), .B2(G283), .ZN(new_n508));
  OR2_X1    g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(KEYINPUT4), .C1(new_n264), .C2(new_n263), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n504), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n267), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n277), .A2(G1), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G257), .A3(new_n270), .ZN(new_n518));
  XNOR2_X1  g0318(.A(KEYINPUT5), .B(G41), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(G274), .A3(new_n270), .A4(new_n514), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(KEYINPUT79), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT79), .B1(new_n518), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n520), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n512), .B2(new_n267), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n524), .A2(G200), .B1(G190), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n521), .B1(new_n267), .B2(new_n512), .ZN(new_n530));
  INV_X1    g0330(.A(new_n525), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n513), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n530), .A2(new_n461), .B1(new_n532), .B2(new_n360), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n495), .A2(new_n497), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n499), .A2(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n271), .A2(G45), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(G250), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n270), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n270), .A2(G274), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(KEYINPUT80), .B1(new_n265), .B2(new_n500), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT81), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n256), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT80), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n259), .A2(new_n548), .A3(G244), .A4(G1698), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n259), .A2(G238), .A3(new_n260), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n541), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n540), .B1(new_n551), .B2(new_n267), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n259), .A2(new_n215), .A3(G68), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n215), .B1(new_n403), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G87), .B2(new_n207), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n298), .B2(new_n485), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n287), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n441), .A2(new_n306), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n496), .A2(new_n441), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n553), .A2(new_n360), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n552), .A2(new_n461), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n496), .A2(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n560), .A3(new_n561), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G190), .B2(new_n552), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n553), .A2(new_n284), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n564), .A2(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n306), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n496), .A2(G107), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n215), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n476), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n546), .A2(new_n215), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n215), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(KEYINPUT22), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n578), .C1(new_n580), .C2(new_n581), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n574), .B1(new_n587), .B2(new_n287), .ZN(new_n588));
  OAI211_X1 g0388(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n259), .A2(KEYINPUT83), .A3(G257), .A4(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n259), .A2(G250), .A3(new_n260), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G33), .A2(G294), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n267), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n517), .A2(G264), .A3(new_n270), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n596), .A2(new_n281), .A3(new_n598), .A4(new_n520), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n539), .A2(new_n517), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n597), .B(new_n600), .C1(new_n595), .C2(new_n267), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n599), .B1(new_n601), .B2(G200), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n588), .A2(new_n602), .A3(KEYINPUT85), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT85), .B1(new_n588), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n535), .B(new_n570), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n587), .A2(new_n287), .ZN(new_n606));
  INV_X1    g0406(.A(new_n574), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n606), .A2(new_n607), .B1(new_n461), .B2(new_n601), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n597), .B1(new_n595), .B2(new_n267), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n520), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n360), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(KEYINPUT84), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n601), .A2(new_n461), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n347), .B1(new_n585), .B2(new_n586), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n574), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT84), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n259), .A2(G257), .A3(new_n260), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n406), .A2(G303), .ZN(new_n620));
  INV_X1    g0420(.A(G264), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n265), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n267), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n517), .A2(new_n270), .ZN(new_n624));
  INV_X1    g0424(.A(G270), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n520), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G169), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n542), .B1(new_n271), .B2(G33), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n393), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(KEYINPUT81), .B(G116), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n292), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n507), .A2(new_n508), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n215), .B1(new_n485), .B2(G33), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n633), .B(new_n287), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n347), .B1(G20), .B2(new_n632), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n640), .B(KEYINPUT20), .C1(new_n635), .C2(new_n636), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n618), .B1(new_n629), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n628), .A2(new_n461), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n634), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n360), .B1(new_n623), .B2(new_n627), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n647), .A2(KEYINPUT21), .A3(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n643), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(G200), .B2(new_n628), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n281), .B2(new_n628), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n612), .A2(new_n617), .A3(new_n651), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n468), .A2(new_n605), .A3(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n317), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n351), .A2(new_n362), .A3(KEYINPUT18), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n368), .B1(new_n367), .B2(new_n361), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n363), .A2(new_n369), .A3(KEYINPUT87), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n429), .A2(new_n460), .A3(new_n462), .A4(new_n452), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n425), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(KEYINPUT88), .ZN(new_n667));
  INV_X1    g0467(.A(new_n378), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n666), .B2(KEYINPUT88), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n664), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n656), .B1(new_n670), .B2(new_n313), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n524), .A2(G179), .B1(G169), .B2(new_n526), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n499), .B1(KEYINPUT86), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT86), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n533), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n673), .A2(new_n570), .A3(new_n674), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n563), .A2(new_n560), .A3(new_n561), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n565), .B(new_n678), .C1(G169), .C2(new_n552), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n552), .A2(G190), .ZN(new_n681));
  INV_X1    g0481(.A(new_n567), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n681), .B(new_n682), .C1(new_n552), .C2(new_n283), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n679), .A2(new_n683), .A3(new_n533), .A4(new_n534), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n680), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n615), .A2(new_n643), .A3(new_n648), .A4(new_n650), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n677), .B(new_n685), .C1(new_n605), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n671), .B1(new_n468), .B2(new_n688), .ZN(G369));
  NAND3_X1  g0489(.A1(new_n271), .A2(new_n215), .A3(G13), .ZN(new_n690));
  OAI21_X1  g0490(.A(G213), .B1(new_n690), .B2(KEYINPUT27), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT27), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n305), .B2(new_n215), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT89), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n305), .A2(new_n692), .A3(new_n215), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT89), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(G213), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(G343), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(G343), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n694), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n647), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n651), .A2(new_n653), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n651), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n615), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n612), .A2(new_n617), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n603), .A2(new_n604), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n588), .A2(new_n703), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n710), .A2(new_n703), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n651), .A2(new_n704), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n712), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n211), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n218), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n687), .A2(new_n730), .A3(new_n703), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n612), .A2(new_n617), .A3(new_n651), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n713), .A3(new_n535), .A4(new_n570), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n679), .B1(new_n684), .B2(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n673), .A2(new_n570), .A3(new_n676), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n734), .B1(KEYINPUT26), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n704), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n731), .B1(new_n737), .B2(new_n730), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  OR3_X1    g0539(.A1(new_n654), .A2(new_n605), .A3(new_n704), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n609), .A2(new_n526), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n644), .A3(KEYINPUT30), .A4(new_n552), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n626), .B1(new_n267), .B2(new_n622), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n552), .A2(new_n745), .A3(G179), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n744), .B1(new_n746), .B2(new_n741), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(G179), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(new_n610), .A3(new_n524), .A4(new_n553), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n704), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n739), .B1(new_n740), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n738), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT92), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n729), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n304), .A2(G20), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n271), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(KEYINPUT93), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n723), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n709), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G330), .B2(new_n707), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n211), .A2(new_n259), .ZN(new_n771));
  INV_X1    g0571(.A(G355), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n211), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n211), .A2(new_n406), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n218), .A2(G45), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n253), .B2(G45), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n773), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n214), .B1(G20), .B2(new_n360), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n768), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(G20), .A2(G179), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n203), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n215), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT32), .ZN(new_n795));
  INV_X1    g0595(.A(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n787), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n790), .B(new_n795), .C1(G68), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G50), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n284), .A2(G190), .A3(new_n791), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT97), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT97), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G87), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n787), .A2(G190), .A3(new_n796), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n319), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n284), .A2(new_n281), .A3(new_n791), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n476), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n281), .A2(G179), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n215), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n485), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n815), .A2(new_n817), .A3(new_n406), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n800), .A2(new_n807), .A3(new_n813), .A4(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n789), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n259), .B(new_n824), .C1(G329), .C2(new_n793), .ZN(new_n825));
  INV_X1    g0625(.A(new_n816), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G283), .A2(new_n826), .B1(new_n799), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(new_n829), .C2(new_n814), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G303), .B2(new_n812), .ZN(new_n831));
  INV_X1    g0631(.A(G326), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n805), .A2(new_n832), .B1(new_n833), .B2(new_n819), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT98), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n822), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n785), .B1(new_n839), .B2(new_n782), .ZN(new_n840));
  INV_X1    g0640(.A(new_n781), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n707), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n770), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  AOI21_X1  g0644(.A(KEYINPUT99), .B1(new_n451), .B2(new_n704), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT99), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n846), .B(new_n703), .C1(new_n446), .C2(new_n450), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n463), .A3(new_n465), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n458), .A2(new_n703), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n452), .A2(new_n460), .A3(new_n462), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(KEYINPUT100), .A3(new_n851), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n688), .B2(new_n704), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n687), .A2(new_n856), .A3(new_n703), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n654), .A2(new_n605), .A3(new_n704), .ZN(new_n861));
  OAI21_X1  g0661(.A(G330), .B1(new_n861), .B2(new_n755), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n768), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n860), .ZN(new_n864));
  INV_X1    g0664(.A(new_n768), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n782), .A2(new_n779), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n203), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n782), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n811), .A2(new_n476), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n259), .B(new_n820), .C1(G311), .C2(new_n793), .ZN(new_n870));
  INV_X1    g0670(.A(new_n814), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G294), .ZN(new_n872));
  INV_X1    g0672(.A(new_n789), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n543), .A2(new_n545), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G283), .A2(new_n799), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n826), .A2(G87), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n870), .A2(new_n872), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n869), .B(new_n877), .C1(G303), .C2(new_n806), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(G143), .ZN(new_n879));
  INV_X1    g0679(.A(G159), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n879), .B1(new_n299), .B2(new_n798), .C1(new_n880), .C2(new_n789), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(G137), .B2(new_n806), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT34), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n826), .A2(G68), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n406), .B1(new_n793), .B2(G132), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(new_n885), .C1(new_n319), .C2(new_n819), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(G50), .B2(new_n812), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n878), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n867), .B1(new_n856), .B2(new_n780), .C1(new_n868), .C2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n864), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(G384));
  OR2_X1    g0691(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(G116), .A4(new_n216), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  NAND4_X1  g0695(.A1(new_n331), .A2(new_n333), .A3(new_n219), .A4(G77), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n202), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n271), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT102), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n660), .A2(new_n668), .A3(new_n662), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n694), .A2(new_n698), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n367), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n367), .A2(new_n361), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n904), .A3(new_n374), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n907), .A2(new_n904), .A3(new_n910), .A4(new_n374), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n348), .A2(new_n349), .B1(new_n289), .B2(new_n290), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n342), .A2(G68), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n335), .A2(new_n337), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n345), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n327), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n374), .B1(new_n918), .B2(new_n362), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n902), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n911), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n920), .B1(new_n370), .B2(new_n378), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n913), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n922), .A2(new_n923), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n925), .B1(new_n930), .B2(new_n924), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n900), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n901), .A2(new_n905), .B1(new_n911), .B2(new_n909), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n925), .B(new_n924), .C1(new_n933), .C2(KEYINPUT38), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT38), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n922), .B2(new_n923), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n934), .B(KEYINPUT102), .C1(new_n925), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT14), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n421), .A3(new_n415), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n395), .A3(new_n703), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n429), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n395), .B(new_n704), .C1(new_n942), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n395), .A2(new_n704), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n425), .A2(new_n429), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n463), .A2(new_n704), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n859), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT101), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n859), .A2(KEYINPUT101), .A3(new_n953), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n930), .A2(new_n924), .ZN(new_n959));
  INV_X1    g0759(.A(new_n664), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n958), .A2(new_n959), .B1(new_n960), .B2(new_n902), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n945), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n738), .A2(new_n467), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n671), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT103), .B1(new_n913), .B2(new_n935), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT103), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n967), .B(new_n924), .C1(new_n933), .C2(KEYINPUT38), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n740), .A2(new_n756), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(KEYINPUT40), .A3(new_n856), .A4(new_n950), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT40), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n950), .B(new_n856), .C1(new_n861), .C2(new_n755), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n937), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n467), .A2(new_n970), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT104), .Z(new_n979));
  AOI21_X1  g0779(.A(new_n739), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n965), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n271), .B2(new_n762), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n965), .A2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n899), .B1(new_n983), .B2(new_n984), .ZN(G367));
  NAND2_X1  g0785(.A1(new_n533), .A2(new_n534), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n673), .A2(new_n676), .A3(new_n704), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n535), .B1(new_n499), .B2(new_n703), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT105), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n986), .B1(new_n991), .B2(new_n712), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n703), .ZN(new_n993));
  INV_X1    g0793(.A(new_n989), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n720), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n682), .A2(new_n703), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  MUX2_X1   g0798(.A(new_n680), .B(new_n570), .S(new_n998), .Z(new_n999));
  AOI22_X1  g0799(.A1(new_n993), .A2(new_n996), .B1(KEYINPUT43), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n991), .A2(new_n717), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT106), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n717), .B2(new_n991), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT106), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1003), .A2(new_n1010), .A3(new_n1006), .A4(new_n1004), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n767), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n758), .B(KEYINPUT92), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n716), .A2(new_n719), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n720), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(KEYINPUT109), .B(new_n708), .C1(new_n1015), .C2(new_n720), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n720), .A2(new_n718), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n989), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT108), .B1(new_n1024), .B2(new_n989), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT108), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1023), .A2(new_n1029), .A3(new_n994), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT44), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n1030), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1027), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n717), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1027), .A2(new_n1033), .A3(new_n717), .A4(new_n1034), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1022), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n760), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n723), .B(KEYINPUT41), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n1013), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1012), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n775), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(new_n246), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n784), .B1(new_n722), .B2(new_n441), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n865), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT46), .B1(new_n812), .B2(new_n874), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G311), .B2(new_n806), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n812), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n259), .B1(new_n793), .B2(G317), .ZN(new_n1051));
  INV_X1    g0851(.A(G283), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n476), .B2(new_n819), .C1(new_n789), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n826), .A2(G97), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n833), .B2(new_n798), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(G303), .C2(new_n871), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1049), .A2(new_n1050), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n816), .A2(new_n203), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n819), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(G68), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n406), .B1(new_n793), .B2(G137), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(new_n798), .C2(new_n880), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1058), .B(new_n1062), .C1(G50), .C2(new_n873), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n806), .A2(G143), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n812), .A2(G58), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n871), .A2(G150), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT47), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n1047), .B1(new_n841), .B2(new_n999), .C1(new_n1069), .C2(new_n868), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT110), .Z(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1043), .A2(new_n1072), .ZN(G387));
  INV_X1    g0873(.A(new_n1021), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n760), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n723), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n716), .A2(new_n841), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n771), .A2(new_n725), .B1(G107), .B2(new_n211), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n242), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1044), .B1(G45), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n725), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT111), .ZN(new_n1083));
  AOI211_X1 g0883(.A(G45), .B(new_n1083), .C1(G68), .C2(G77), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n323), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT50), .B1(new_n323), .B2(new_n202), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1084), .B1(KEYINPUT111), .B2(new_n1082), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1079), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n768), .B1(new_n1088), .B2(new_n784), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G68), .A2(new_n873), .B1(new_n799), .B2(new_n323), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1059), .A2(new_n441), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n406), .B1(new_n793), .B2(G150), .ZN(new_n1092));
  AND4_X1   g0892(.A1(new_n1054), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n806), .A2(G159), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n812), .A2(G77), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n871), .A2(G50), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n871), .A2(G317), .B1(new_n873), .B2(G303), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT112), .Z(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n823), .B2(new_n798), .C1(new_n829), .C2(new_n805), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT48), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n811), .A2(new_n833), .B1(new_n1052), .B2(new_n819), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1102), .A2(KEYINPUT49), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n259), .B1(new_n793), .B2(G326), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(new_n632), .C2(new_n816), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT49), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1097), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1089), .B1(new_n1109), .B2(new_n782), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1074), .A2(new_n767), .B1(new_n1078), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1077), .A2(new_n1111), .ZN(G393));
  NAND3_X1  g0912(.A1(new_n1037), .A2(KEYINPUT113), .A3(new_n1038), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1035), .A2(new_n1114), .A3(new_n1036), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1039), .B(new_n723), .C1(new_n1116), .C2(new_n1022), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G50), .A2(new_n799), .B1(new_n873), .B2(new_n323), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1059), .A2(G77), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n406), .B1(new_n793), .B2(G143), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1118), .A2(new_n876), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n805), .A2(new_n299), .B1(new_n880), .B2(new_n814), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT51), .Z(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(new_n221), .C2(new_n812), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n806), .A2(G317), .B1(G311), .B2(new_n871), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n406), .B1(new_n792), .B2(new_n829), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1127), .B(new_n817), .C1(new_n874), .C2(new_n1059), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G294), .A2(new_n873), .B1(new_n799), .B2(G303), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n1052), .C2(new_n811), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n782), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n775), .A2(new_n250), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n783), .C1(new_n485), .C2(new_n211), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n768), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n781), .B2(new_n991), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n1116), .B2(new_n767), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1117), .A2(new_n1137), .ZN(G390));
  OAI211_X1 g0938(.A(new_n932), .B(new_n938), .C1(new_n958), .C2(new_n944), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n970), .A2(G330), .A3(new_n856), .A4(new_n950), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n952), .B1(new_n737), .B2(new_n856), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n969), .B(new_n943), .C1(new_n951), .C2(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n951), .B1(new_n862), .B2(new_n857), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n1140), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n956), .A2(new_n957), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n757), .A2(KEYINPUT114), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT114), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n857), .B1(new_n862), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n950), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n757), .A2(new_n467), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n671), .A2(new_n963), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g0958(.A1(new_n1143), .A2(new_n1144), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n724), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1140), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT115), .B1(new_n1165), .B2(new_n1158), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT115), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n951), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1153), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1156), .B1(new_n1171), .B2(new_n1148), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1167), .B(new_n1172), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1160), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1165), .A2(new_n1013), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n866), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n873), .A2(G97), .B1(G77), .B2(new_n1059), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n476), .B2(new_n798), .C1(new_n542), .C2(new_n814), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n884), .B1(new_n833), .B2(new_n792), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT118), .Z(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(G283), .C2(new_n806), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n813), .A2(new_n406), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT117), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n812), .A2(G150), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G132), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n814), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n406), .B1(new_n793), .B2(G125), .ZN(new_n1189));
  INV_X1    g0989(.A(G137), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1189), .B1(new_n880), .B2(new_n819), .C1(new_n798), .C2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n816), .A2(new_n202), .B1(new_n789), .B2(new_n1192), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1186), .A2(new_n1188), .A3(new_n1191), .A4(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1184), .A2(new_n1185), .B1(new_n806), .B2(G128), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1181), .A2(new_n1183), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n768), .B1(new_n323), .B2(new_n1176), .C1(new_n1196), .C2(new_n868), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n939), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n779), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1175), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1174), .A2(new_n1200), .ZN(G378));
  XOR2_X1   g1001(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n307), .A2(new_n903), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT120), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n313), .A2(new_n317), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1205), .B1(new_n313), .B2(new_n317), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1203), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1202), .A3(new_n1206), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n976), .A2(G330), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n973), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n971), .B1(new_n966), .B2(new_n968), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n976), .A2(G330), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1212), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n958), .A2(new_n959), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n960), .A2(new_n902), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n943), .B1(new_n932), .B2(new_n938), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1214), .A2(new_n1218), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n973), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n945), .A3(new_n1225), .A4(new_n961), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1013), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1217), .A2(new_n779), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n768), .B1(G50), .B2(new_n1176), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n259), .A2(G41), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G50), .B(new_n1230), .C1(new_n256), .C2(new_n276), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n826), .A2(G58), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n485), .B2(new_n798), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1060), .B(new_n1230), .C1(new_n1052), .C2(new_n792), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n873), .B2(new_n441), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(G107), .C2(new_n871), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n1095), .C1(new_n542), .C2(new_n805), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT58), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n806), .A2(G125), .B1(G150), .B2(new_n1059), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT119), .Z(new_n1242));
  OAI22_X1  g1042(.A1(new_n1187), .A2(new_n798), .B1(new_n789), .B2(new_n1190), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G128), .B2(new_n871), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n811), .C2(new_n1192), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT59), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n880), .B2(new_n816), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1240), .B1(new_n1239), .B2(new_n1238), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1229), .B1(new_n1249), .B2(new_n782), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1227), .B1(new_n1228), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT57), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1159), .B2(new_n1156), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT121), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1253), .B(KEYINPUT121), .C1(new_n1159), .C2(new_n1156), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1163), .A2(new_n1164), .A3(new_n1172), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1259), .A2(new_n1157), .B1(new_n1226), .B2(new_n1223), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n723), .B1(new_n1260), .B2(KEYINPUT57), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1251), .B1(new_n1258), .B2(new_n1261), .ZN(G375));
  NAND3_X1  g1062(.A1(new_n1171), .A2(new_n1148), .A3(new_n1156), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1041), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1158), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n951), .A2(new_n779), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n768), .B1(G68), .B2(new_n1176), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n259), .B1(new_n793), .B2(G303), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1091), .A2(new_n1268), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n476), .A2(new_n789), .B1(new_n798), .B2(new_n632), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1058), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n485), .B2(new_n811), .C1(new_n1052), .C2(new_n814), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n805), .A2(new_n833), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n789), .A2(new_n299), .B1(new_n202), .B2(new_n819), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT122), .Z(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n880), .B2(new_n811), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n798), .A2(new_n1192), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n406), .B1(new_n793), .B2(G128), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1232), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n1190), .B2(new_n814), .C1(new_n1187), .C2(new_n805), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1272), .A2(new_n1273), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1267), .B1(new_n1281), .B2(new_n782), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1154), .A2(new_n767), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1265), .A2(new_n1283), .ZN(G381));
  OR2_X1    g1084(.A1(G375), .A2(G378), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1077), .A2(new_n843), .A3(new_n1111), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n890), .ZN(new_n1287));
  OR3_X1    g1087(.A1(G390), .A2(new_n1287), .A3(G381), .ZN(new_n1288));
  OR3_X1    g1088(.A1(new_n1285), .A2(G387), .A3(new_n1288), .ZN(G407));
  NAND3_X1  g1089(.A1(new_n700), .A2(new_n701), .A3(G213), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G407), .B(G213), .C1(new_n1285), .C2(new_n1290), .ZN(G409));
  AOI21_X1  g1091(.A(new_n843), .B1(new_n1077), .B2(new_n1111), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(G390), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1117), .B(new_n1137), .C1(new_n1286), .C2(new_n1292), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(G387), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1294), .A2(new_n1043), .A3(new_n1072), .A4(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1251), .C1(new_n1258), .C2(new_n1261), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1251), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1174), .A3(new_n1200), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1290), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1290), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1154), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1307), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1156), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n1148), .A4(new_n1156), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT123), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1263), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n724), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1308), .A2(new_n1311), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1315), .A2(G384), .A3(new_n1283), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G384), .B1(new_n1315), .B2(new_n1283), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G2897), .B(new_n1306), .C1(new_n1318), .C2(KEYINPUT124), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT124), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1306), .A2(G2897), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1320), .B(new_n1321), .C1(new_n1316), .C2(new_n1317), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1319), .A2(new_n1322), .B1(KEYINPUT124), .B2(new_n1318), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1305), .B2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1304), .A2(new_n1290), .A3(new_n1318), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1299), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT125), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1315), .A2(new_n1283), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n890), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1315), .A2(G384), .A3(new_n1283), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1304), .A2(new_n1290), .A3(new_n1336), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1306), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1318), .A2(KEYINPUT124), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1321), .B1(new_n1334), .B2(new_n1320), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1322), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1342), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1340), .B1(new_n1341), .B2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1339), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1325), .A2(new_n1335), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1330), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1299), .B1(new_n1341), .B2(new_n1336), .ZN(new_n1350));
  AND4_X1   g1150(.A1(new_n1330), .A2(new_n1324), .A3(new_n1350), .A4(new_n1348), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1329), .B1(new_n1349), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(KEYINPUT126), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1354), .B(new_n1329), .C1(new_n1349), .C2(new_n1351), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(G405));
  NAND3_X1  g1156(.A1(G375), .A2(new_n1174), .A3(new_n1200), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1300), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1318), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1357), .A2(new_n1300), .A3(new_n1334), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1359), .A2(new_n1299), .A3(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1299), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT127), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1361), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1364), .B1(new_n1363), .B2(new_n1362), .ZN(G402));
endmodule


