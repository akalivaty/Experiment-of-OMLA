

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n405) );
  XNOR2_X1 U323 ( .A(n467), .B(KEYINPUT94), .ZN(n482) );
  XOR2_X1 U324 ( .A(n398), .B(n397), .Z(n567) );
  XOR2_X1 U325 ( .A(n462), .B(KEYINPUT28), .Z(n521) );
  XNOR2_X1 U326 ( .A(n419), .B(n418), .ZN(n509) );
  XOR2_X1 U327 ( .A(KEYINPUT80), .B(KEYINPUT17), .Z(n290) );
  AND2_X1 U328 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  INV_X1 U329 ( .A(KEYINPUT25), .ZN(n453) );
  XNOR2_X1 U330 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n422) );
  XNOR2_X1 U331 ( .A(n423), .B(n422), .ZN(n441) );
  XNOR2_X1 U332 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U333 ( .A(n413), .B(n291), .ZN(n414) );
  XNOR2_X1 U334 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U335 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U336 ( .A(n377), .B(n376), .ZN(n380) );
  XNOR2_X1 U337 ( .A(KEYINPUT38), .B(n485), .ZN(n492) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n444) );
  XNOR2_X1 U339 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n293) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G85GAT), .ZN(n350) );
  INV_X1 U342 ( .A(n350), .ZN(n292) );
  XOR2_X1 U343 ( .A(n293), .B(n292), .Z(n307) );
  XNOR2_X1 U344 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n294), .B(G162GAT), .ZN(n343) );
  XOR2_X1 U346 ( .A(G106GAT), .B(n343), .Z(n296) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U349 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n298) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G43GAT), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n390) );
  XNOR2_X1 U356 ( .A(G36GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n303), .B(G218GAT), .ZN(n409) );
  XNOR2_X1 U358 ( .A(n390), .B(n409), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U360 ( .A(n307), .B(n306), .Z(n533) );
  XOR2_X1 U361 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n309) );
  XNOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U364 ( .A(n310), .B(G127GAT), .Z(n312) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G120GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n427) );
  XOR2_X1 U367 ( .A(G183GAT), .B(G99GAT), .Z(n314) );
  XNOR2_X1 U368 ( .A(G43GAT), .B(G190GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U370 ( .A(KEYINPUT79), .B(G71GAT), .Z(n316) );
  XNOR2_X1 U371 ( .A(G15GAT), .B(G176GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U373 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U374 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n320) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U377 ( .A(KEYINPUT20), .B(n321), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n427), .B(n324), .ZN(n328) );
  XNOR2_X1 U380 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n290), .B(n325), .ZN(n326) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(n326), .ZN(n410) );
  INV_X1 U383 ( .A(n410), .ZN(n327) );
  XOR2_X2 U384 ( .A(n328), .B(n327), .Z(n523) );
  XOR2_X1 U385 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n330) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n430) );
  XOR2_X1 U388 ( .A(G78GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U389 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U390 ( .A(n332), .B(n331), .ZN(n355) );
  XNOR2_X1 U391 ( .A(n430), .B(n355), .ZN(n347) );
  XOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .Z(n364) );
  XOR2_X1 U393 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n334) );
  XNOR2_X1 U394 ( .A(G218GAT), .B(KEYINPUT85), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U396 ( .A(n364), .B(n335), .Z(n337) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U399 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n339) );
  XNOR2_X1 U400 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U402 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n342), .B(G211GAT), .ZN(n418) );
  XNOR2_X1 U405 ( .A(n343), .B(n418), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n462) );
  XOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT32), .Z(n349) );
  XNOR2_X1 U409 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n353) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n354), .B(KEYINPUT70), .ZN(n357) );
  XOR2_X1 U415 ( .A(n355), .B(KEYINPUT33), .Z(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n363) );
  XOR2_X1 U417 ( .A(G57GAT), .B(KEYINPUT67), .Z(n359) );
  XNOR2_X1 U418 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n378) );
  XOR2_X1 U420 ( .A(G64GAT), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(G204GAT), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n417) );
  XOR2_X1 U423 ( .A(n378), .B(n417), .Z(n362) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n448) );
  INV_X1 U425 ( .A(n448), .ZN(n572) );
  XOR2_X1 U426 ( .A(G8GAT), .B(G183GAT), .Z(n413) );
  XOR2_X1 U427 ( .A(n413), .B(n364), .Z(n366) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n368) );
  XNOR2_X1 U431 ( .A(G64GAT), .B(KEYINPUT73), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n377) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G1GAT), .Z(n393) );
  XOR2_X1 U435 ( .A(KEYINPUT75), .B(G78GAT), .Z(n372) );
  XNOR2_X1 U436 ( .A(G127GAT), .B(G211GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U438 ( .A(n393), .B(n373), .Z(n375) );
  INV_X1 U439 ( .A(KEYINPUT12), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n378), .B(KEYINPUT15), .ZN(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n577) );
  INV_X1 U442 ( .A(n577), .ZN(n548) );
  XOR2_X1 U443 ( .A(KEYINPUT36), .B(n533), .Z(n582) );
  NOR2_X1 U444 ( .A1(n548), .A2(n582), .ZN(n381) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n381), .Z(n382) );
  XNOR2_X1 U446 ( .A(n382), .B(KEYINPUT64), .ZN(n383) );
  NOR2_X1 U447 ( .A1(n572), .A2(n383), .ZN(n399) );
  XOR2_X1 U448 ( .A(G197GAT), .B(G22GAT), .Z(n385) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(G113GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U451 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n387) );
  XNOR2_X1 U452 ( .A(G141GAT), .B(G8GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT29), .ZN(n392) );
  NAND2_X1 U456 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n396) );
  XNOR2_X1 U459 ( .A(G50GAT), .B(G36GAT), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  INV_X1 U461 ( .A(n567), .ZN(n540) );
  NAND2_X1 U462 ( .A1(n399), .A2(n540), .ZN(n408) );
  XOR2_X1 U463 ( .A(n572), .B(KEYINPUT41), .Z(n557) );
  NAND2_X1 U464 ( .A1(n557), .A2(n567), .ZN(n401) );
  XOR2_X1 U465 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U467 ( .A(n577), .B(KEYINPUT107), .Z(n561) );
  NOR2_X1 U468 ( .A1(n402), .A2(n561), .ZN(n403) );
  XNOR2_X1 U469 ( .A(n403), .B(KEYINPUT109), .ZN(n404) );
  NOR2_X1 U470 ( .A1(n533), .A2(n404), .ZN(n406) );
  NAND2_X1 U471 ( .A1(n408), .A2(n407), .ZN(n518) );
  XNOR2_X1 U472 ( .A(n518), .B(KEYINPUT48), .ZN(n421) );
  XOR2_X1 U473 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n412) );
  XOR2_X1 U474 ( .A(n410), .B(n409), .Z(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U477 ( .A(KEYINPUT118), .B(n509), .Z(n420) );
  NAND2_X1 U478 ( .A1(n421), .A2(n420), .ZN(n423) );
  XOR2_X1 U479 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n425) );
  XNOR2_X1 U480 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n440) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G155GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n438) );
  XOR2_X1 U486 ( .A(KEYINPUT87), .B(n430), .Z(n432) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U489 ( .A(KEYINPUT6), .B(G57GAT), .Z(n434) );
  XNOR2_X1 U490 ( .A(G1GAT), .B(G148GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U492 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n458) );
  INV_X1 U495 ( .A(n458), .ZN(n505) );
  NAND2_X1 U496 ( .A1(n441), .A2(n505), .ZN(n565) );
  NOR2_X1 U497 ( .A1(n462), .A2(n565), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n442), .B(KEYINPUT55), .ZN(n443) );
  NOR2_X2 U499 ( .A1(n523), .A2(n443), .ZN(n560) );
  NAND2_X1 U500 ( .A1(n533), .A2(n560), .ZN(n445) );
  XOR2_X1 U501 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n447) );
  XNOR2_X1 U502 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n472) );
  NAND2_X1 U504 ( .A1(n567), .A2(n448), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n449), .B(KEYINPUT71), .ZN(n484) );
  NAND2_X1 U506 ( .A1(n523), .A2(n462), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n450), .B(KEYINPUT92), .ZN(n451) );
  XOR2_X1 U508 ( .A(KEYINPUT26), .B(n451), .Z(n539) );
  INV_X1 U509 ( .A(n539), .ZN(n564) );
  XNOR2_X1 U510 ( .A(KEYINPUT27), .B(n509), .ZN(n460) );
  NOR2_X1 U511 ( .A1(n564), .A2(n460), .ZN(n456) );
  NOR2_X1 U512 ( .A1(n509), .A2(n523), .ZN(n452) );
  NOR2_X1 U513 ( .A1(n462), .A2(n452), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT93), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n460), .A2(n505), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT91), .ZN(n519) );
  INV_X1 U520 ( .A(n521), .ZN(n463) );
  NOR2_X1 U521 ( .A1(n519), .A2(n463), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n464), .A2(n523), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n469) );
  INV_X1 U525 ( .A(n533), .ZN(n551) );
  NAND2_X1 U526 ( .A1(n551), .A2(n577), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  AND2_X1 U528 ( .A1(n482), .A2(n470), .ZN(n494) );
  NAND2_X1 U529 ( .A1(n484), .A2(n494), .ZN(n478) );
  NOR2_X1 U530 ( .A1(n505), .A2(n478), .ZN(n471) );
  XOR2_X1 U531 ( .A(n472), .B(n471), .Z(G1324GAT) );
  NOR2_X1 U532 ( .A1(n509), .A2(n478), .ZN(n474) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(G1325GAT) );
  NOR2_X1 U535 ( .A1(n523), .A2(n478), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT35), .B(KEYINPUT98), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(G15GAT), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U539 ( .A1(n521), .A2(n478), .ZN(n480) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1327GAT) );
  NOR2_X1 U542 ( .A1(n582), .A2(n577), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n483), .ZN(n504) );
  NAND2_X1 U545 ( .A1(n504), .A2(n484), .ZN(n485) );
  NOR2_X1 U546 ( .A1(n492), .A2(n505), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n509), .A2(n492), .ZN(n488) );
  XOR2_X1 U550 ( .A(G36GAT), .B(n488), .Z(G1329GAT) );
  NOR2_X1 U551 ( .A1(n492), .A2(n523), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U554 ( .A(G43GAT), .B(n491), .Z(G1330GAT) );
  NOR2_X1 U555 ( .A1(n521), .A2(n492), .ZN(n493) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n493), .Z(G1331GAT) );
  INV_X1 U557 ( .A(n557), .ZN(n543) );
  NOR2_X1 U558 ( .A1(n543), .A2(n567), .ZN(n503) );
  NAND2_X1 U559 ( .A1(n503), .A2(n494), .ZN(n500) );
  NOR2_X1 U560 ( .A1(n505), .A2(n500), .ZN(n496) );
  XNOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT42), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n497), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n509), .A2(n500), .ZN(n498) );
  XOR2_X1 U565 ( .A(G64GAT), .B(n498), .Z(G1333GAT) );
  NOR2_X1 U566 ( .A1(n523), .A2(n500), .ZN(n499) );
  XOR2_X1 U567 ( .A(G71GAT), .B(n499), .Z(G1334GAT) );
  NOR2_X1 U568 ( .A1(n521), .A2(n500), .ZN(n502) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n504), .A2(n503), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n505), .A2(n514), .ZN(n507) );
  XNOR2_X1 U573 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n509), .A2(n514), .ZN(n510) );
  XOR2_X1 U577 ( .A(KEYINPUT104), .B(n510), .Z(n511) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n511), .ZN(G1337GAT) );
  NOR2_X1 U579 ( .A1(n523), .A2(n514), .ZN(n513) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT105), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(G1338GAT) );
  NOR2_X1 U582 ( .A1(n521), .A2(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(KEYINPUT106), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n517), .Z(G1339GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n525) );
  XOR2_X1 U587 ( .A(n518), .B(KEYINPUT48), .Z(n520) );
  NOR2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n538) );
  NAND2_X1 U589 ( .A1(n521), .A2(n538), .ZN(n522) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n534), .A2(n567), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U595 ( .A1(n534), .A2(n557), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n531) );
  NAND2_X1 U599 ( .A1(n534), .A2(n561), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U603 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n537), .Z(G1343GAT) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n540), .A2(n550), .ZN(n541) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n541), .Z(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT116), .B(n542), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n550), .A2(n543), .ZN(n547) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n550), .ZN(n549) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  NAND2_X1 U619 ( .A1(n567), .A2(n560), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT123), .B(n566), .ZN(n581) );
  INV_X1 U632 ( .A(n581), .ZN(n578) );
  NAND2_X1 U633 ( .A1(n567), .A2(n578), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U639 ( .A1(n578), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

