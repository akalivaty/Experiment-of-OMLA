//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n534, new_n535,
    new_n536, new_n537, new_n539, new_n540, new_n542, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  AOI22_X1  g034(.A1(G567), .A2(new_n458), .B1(new_n459), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n464), .B2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n462), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(new_n472), .A3(new_n461), .A4(new_n465), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g052(.A(KEYINPUT69), .B(new_n469), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n471), .A2(new_n472), .A3(G2105), .A4(new_n465), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n481), .B1(new_n473), .B2(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  OR2_X1    g062(.A1(KEYINPUT70), .A2(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT70), .A2(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n461), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n484), .A2(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n473), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n463), .A2(new_n465), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n494), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n502), .A2(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(G88), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n511), .A2(G89), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(G168));
  AOI22_X1  g098(.A1(new_n511), .A2(G90), .B1(new_n513), .B2(G52), .ZN(new_n524));
  INV_X1    g099(.A(G64), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n502), .B2(new_n504), .ZN(new_n526));
  AND2_X1   g101(.A1(G77), .A2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n524), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n511), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n507), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT74), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT75), .Z(G176));
  XOR2_X1   g116(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n542));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n539), .A2(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n511), .A2(G91), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n513), .A2(G53), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(KEYINPUT9), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(KEYINPUT9), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n546), .B1(new_n507), .B2(new_n547), .C1(new_n549), .C2(new_n550), .ZN(G299));
  INV_X1    g126(.A(new_n532), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n531), .B1(new_n524), .B2(new_n528), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n554));
  NOR3_X1   g129(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT77), .B1(new_n530), .B2(new_n532), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  NAND2_X1  g133(.A1(new_n511), .A2(G87), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n513), .A2(G49), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(new_n505), .A2(G61), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT78), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n511), .A2(G86), .B1(new_n513), .B2(G48), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G305));
  AOI22_X1  g144(.A1(new_n511), .A2(G85), .B1(new_n513), .B2(G47), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT80), .Z(new_n571));
  AOI22_X1  g146(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n507), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(new_n505), .A2(G66), .ZN(new_n576));
  INV_X1    g151(.A(G79), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n501), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n579));
  INV_X1    g154(.A(new_n511), .ZN(new_n580));
  INV_X1    g155(.A(G92), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(G301), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(G868), .ZN(G321));
  XOR2_X1   g164(.A(G321), .B(KEYINPUT82), .Z(G284));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(G299), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n591), .B2(G168), .ZN(G297));
  OAI21_X1  g168(.A(new_n592), .B1(new_n591), .B2(G168), .ZN(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n585), .B1(new_n595), .B2(G860), .ZN(G148));
  INV_X1    g171(.A(new_n537), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(new_n591), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n586), .A2(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n591), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n496), .A2(G2104), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT13), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(G2100), .ZN(new_n605));
  INV_X1    g180(.A(new_n473), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G135), .ZN(new_n607));
  INV_X1    g182(.A(new_n484), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G123), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n461), .A2(KEYINPUT83), .A3(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT83), .B1(new_n461), .B2(G111), .ZN(new_n611));
  OR2_X1    g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(G2104), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n607), .B(new_n609), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n605), .A2(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(G2427), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2430), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(KEYINPUT14), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(G1341), .B(G1348), .Z(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2451), .B(G2454), .Z(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n629), .ZN(new_n631));
  AND3_X1   g206(.A1(new_n630), .A2(G14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT85), .Z(G401));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n634), .B1(new_n636), .B2(KEYINPUT87), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(KEYINPUT87), .B2(new_n636), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT88), .B(KEYINPUT17), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n635), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n634), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n638), .B(new_n640), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n639), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n636), .A2(new_n634), .A3(new_n639), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n644), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2096), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  AND2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n654), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G229));
  NAND2_X1  g244(.A1(new_n585), .A2(G16), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(G4), .B2(G16), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT95), .B(G1348), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT24), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n675), .B2(G34), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n675), .B2(G34), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G160), .B2(G29), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(G2084), .ZN(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NOR2_X1   g255(.A1(G286), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT101), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g258(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G1966), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n674), .A2(G26), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT98), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  OR2_X1    g264(.A1(G104), .A2(G2105), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n690), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n691));
  INV_X1    g266(.A(G128), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n484), .B2(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n606), .B2(G140), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n694), .B2(new_n674), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT99), .B(G2067), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n673), .A2(new_n679), .A3(new_n686), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n685), .A2(G1966), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n606), .A2(G139), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT25), .Z(new_n702));
  INV_X1    g277(.A(new_n495), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n703), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n700), .B(new_n702), .C1(new_n461), .C2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G33), .B(new_n705), .S(G29), .Z(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G2072), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT30), .B(G28), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n708), .A2(new_n674), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n614), .B2(new_n674), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n706), .B2(G2072), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n671), .A2(new_n672), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n699), .A2(new_n707), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT91), .B(G16), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G20), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT23), .Z(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G299), .B2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G1956), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n674), .A2(G32), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT100), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT26), .ZN(new_n725));
  AOI22_X1  g300(.A1(G141), .A2(new_n606), .B1(new_n608), .B2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(new_n674), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n698), .A2(new_n715), .A3(new_n721), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n674), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n674), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT104), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT103), .B(G2078), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n716), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n537), .B2(new_n738), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT96), .B(G1341), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT97), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT105), .B(KEYINPUT29), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n743), .B(new_n749), .C1(G2084), .C2(new_n678), .ZN(new_n750));
  NOR2_X1   g325(.A1(G5), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G171), .B2(G16), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT102), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n732), .A2(new_n737), .A3(new_n750), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n680), .A2(G6), .ZN(new_n757));
  INV_X1    g332(.A(G305), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(new_n680), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  XOR2_X1   g335(.A(KEYINPUT32), .B(G1981), .Z(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n716), .A2(G22), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT93), .Z(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G303), .B2(new_n738), .ZN(new_n765));
  INV_X1    g340(.A(G1971), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n680), .A2(G23), .ZN(new_n769));
  INV_X1    g344(.A(G288), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n680), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT33), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1976), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n760), .A2(new_n761), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n768), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT34), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  MUX2_X1   g353(.A(G24), .B(G290), .S(new_n738), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1986), .ZN(new_n780));
  NOR2_X1   g355(.A1(G25), .A2(G29), .ZN(new_n781));
  OAI21_X1  g356(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n784));
  OAI221_X1 g359(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G119), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n484), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G131), .B2(new_n606), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n781), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n780), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n777), .A2(new_n778), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT36), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n797), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n756), .B1(new_n798), .B2(new_n799), .ZN(G311));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  INV_X1    g376(.A(new_n756), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(G150));
  NAND2_X1  g378(.A1(new_n513), .A2(G55), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT106), .B(G93), .Z(new_n805));
  AOI22_X1  g380(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n804), .B1(new_n580), .B2(new_n805), .C1(new_n806), .C2(new_n507), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n536), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n597), .B2(new_n807), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n586), .A2(new_n595), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n813));
  AOI21_X1  g388(.A(G860), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n807), .A2(G860), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT107), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT37), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(G145));
  INV_X1    g394(.A(new_n694), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n705), .A2(KEYINPUT108), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n728), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n494), .A2(new_n498), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT70), .B(G114), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n491), .B1(new_n824), .B2(G2105), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n608), .B2(G126), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n728), .A2(new_n821), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n822), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n827), .B1(new_n822), .B2(new_n828), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n608), .A2(G130), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n461), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G142), .B2(new_n606), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n603), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n788), .ZN(new_n839));
  INV_X1    g414(.A(new_n831), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n840), .A2(new_n694), .A3(new_n829), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n832), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT109), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n832), .A2(new_n841), .ZN(new_n844));
  INV_X1    g419(.A(new_n839), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(KEYINPUT109), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G160), .B(new_n485), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n614), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT110), .B(G37), .Z(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n844), .B2(new_n845), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n842), .A2(KEYINPUT111), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT111), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n839), .A2(new_n832), .A3(new_n841), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT112), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT112), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n851), .B(new_n852), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT113), .B(KEYINPUT40), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(G395));
  XOR2_X1   g437(.A(new_n809), .B(new_n599), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n585), .B(G299), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT41), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT42), .ZN(new_n868));
  XNOR2_X1  g443(.A(G290), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(G303), .B(new_n770), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT42), .B1(new_n866), .B2(new_n867), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n868), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n868), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(G868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n807), .A2(new_n591), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(G295));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n876), .ZN(G331));
  INV_X1    g453(.A(new_n871), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT116), .ZN(new_n880));
  NOR2_X1   g455(.A1(G171), .A2(G168), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT114), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n882), .B(new_n883), .C1(G301), .C2(G286), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n554), .B1(new_n552), .B2(new_n553), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n530), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n886));
  AOI21_X1  g461(.A(G286), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT114), .B1(new_n887), .B2(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n888), .A3(new_n809), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(new_n864), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n888), .ZN(new_n891));
  INV_X1    g466(.A(new_n809), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n880), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n864), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n809), .B1(new_n884), .B2(new_n888), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n895), .A2(KEYINPUT116), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT115), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(KEYINPUT115), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n889), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n865), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n879), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n890), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n893), .A2(new_n889), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n879), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n852), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n905), .A2(new_n906), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n909), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n871), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT43), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n905), .A2(KEYINPUT43), .A3(new_n911), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n906), .B1(new_n914), .B2(new_n916), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(G397));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G164), .B2(G1384), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n477), .A2(new_n478), .ZN(new_n926));
  INV_X1    g501(.A(new_n468), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT117), .B(G40), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n728), .B(G1996), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n694), .B(G2067), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n788), .A2(new_n790), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n788), .A2(new_n790), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G290), .B(G1986), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT54), .ZN(new_n939));
  INV_X1    g514(.A(G2078), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n827), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n930), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n823), .B2(new_n826), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT45), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT118), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n468), .B(new_n928), .C1(new_n477), .C2(new_n478), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n945), .A2(new_n925), .A3(new_n947), .A4(KEYINPUT118), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n940), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(KEYINPUT126), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT126), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT118), .ZN(new_n954));
  OAI211_X1 g529(.A(G160), .B(new_n929), .C1(new_n944), .C2(KEYINPUT45), .ZN(new_n955));
  NOR3_X1   g530(.A1(G164), .A2(new_n924), .A3(G1384), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G2078), .B1(new_n957), .B2(new_n948), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n958), .B2(KEYINPUT53), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n945), .A2(new_n925), .A3(new_n947), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(KEYINPUT53), .A3(new_n940), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n472), .A2(new_n465), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(G138), .A3(new_n461), .A4(new_n471), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n965), .A2(KEYINPUT4), .B1(new_n496), .B2(new_n497), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n963), .B(new_n941), .C1(new_n966), .C2(new_n492), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT119), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n944), .A2(KEYINPUT119), .A3(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n827), .A2(new_n941), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n930), .B1(KEYINPUT50), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n754), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n952), .A2(new_n959), .A3(new_n962), .A4(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n976), .A2(new_n588), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n940), .A2(KEYINPUT53), .A3(G40), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n945), .A2(new_n925), .A3(G160), .A4(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n952), .A2(new_n959), .A3(new_n975), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(new_n588), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n939), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n957), .A2(new_n766), .A3(new_n948), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n973), .A2(new_n748), .A3(new_n967), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(G8), .B1(new_n930), .B2(new_n972), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT120), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT120), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(G8), .C1(new_n930), .C2(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G305), .A2(G1981), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n567), .A2(new_n996), .A3(new_n568), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT49), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n994), .A2(new_n999), .A3(KEYINPUT121), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n985), .B1(G2090), .B2(new_n974), .ZN(new_n1005));
  INV_X1    g580(.A(new_n984), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(G8), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n770), .A2(G1976), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n994), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n770), .B2(G1976), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1009), .B(new_n1012), .C1(new_n991), .C2(new_n993), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n989), .A2(new_n1004), .A3(new_n1007), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1348), .B1(new_n971), .B2(new_n973), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n586), .A2(KEYINPUT60), .ZN(new_n1017));
  INV_X1    g592(.A(G2067), .ZN(new_n1018));
  NAND4_X1  g593(.A1(G160), .A2(new_n944), .A3(new_n1018), .A4(new_n929), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n947), .A2(KEYINPUT122), .A3(new_n1018), .A4(new_n944), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1016), .A2(new_n1017), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G299), .B(KEYINPUT57), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1956), .B1(new_n973), .B2(new_n967), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n960), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1025), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n947), .A3(new_n967), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n720), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G299), .B(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1033), .B(new_n1035), .C1(new_n960), .C2(new_n1028), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1024), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n961), .A2(new_n1027), .B1(new_n1032), .B2(new_n720), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(new_n1035), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1025), .A2(KEYINPUT123), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1042), .B(new_n1044), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT58), .B(G1341), .Z(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n930), .B2(new_n972), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n960), .B2(G1996), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n537), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT59), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(new_n1051), .A3(new_n537), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1041), .A2(new_n1045), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1348), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n974), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1023), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n586), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1016), .A2(new_n585), .A3(new_n1023), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT60), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1039), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1045), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1036), .B1(new_n1061), .B2(new_n1057), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1015), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G2084), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n971), .A2(new_n973), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1966), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n960), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(G168), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT125), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1068), .A2(new_n1073), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT124), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1069), .A2(new_n1076), .A3(new_n1070), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n988), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(G286), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n980), .A2(G171), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(KEYINPUT54), .C1(new_n588), .C2(new_n976), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n982), .A2(new_n1063), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G288), .A2(G1976), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1004), .A2(new_n1085), .B1(new_n996), .B2(new_n758), .ZN(new_n1086));
  INV_X1    g661(.A(new_n994), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1004), .A2(new_n1014), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1086), .A2(new_n1087), .B1(new_n1007), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1079), .A2(G168), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1015), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1004), .A2(new_n1007), .A3(new_n1014), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1006), .B1(new_n1005), .B2(G8), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1089), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1084), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1078), .A2(new_n1099), .A3(new_n1080), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n977), .A2(new_n1093), .A3(new_n989), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n938), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n931), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(G1996), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT46), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n933), .A2(new_n728), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1106), .A2(new_n1107), .B1(new_n931), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT47), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n932), .A2(new_n788), .A3(new_n790), .A4(new_n933), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n694), .A2(new_n1018), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1105), .A2(G1986), .A3(G290), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n936), .A2(new_n931), .B1(new_n1115), .B2(KEYINPUT48), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1115), .A2(KEYINPUT48), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT127), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1104), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g696(.A1(new_n651), .A2(G319), .ZN(new_n1123));
  NOR3_X1   g697(.A1(G229), .A2(new_n632), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g698(.A(new_n860), .B(new_n1124), .C1(new_n920), .C2(new_n921), .ZN(G225));
  INV_X1    g699(.A(G225), .ZN(G308));
endmodule


