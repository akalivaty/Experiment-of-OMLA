//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n449, new_n451, new_n455,
    new_n456, new_n457, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  NAND2_X1  g023(.A1(G94), .A2(G452), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(G160));
  NOR2_X1   g052(.A1(new_n463), .A2(new_n464), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(G162));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n463), .B2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n489), .B(new_n492), .C1(new_n464), .C2(new_n463), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT70), .A2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT70), .A2(G114), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n495), .B(G2105), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(KEYINPUT70), .A2(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n462), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G102), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT71), .B1(new_n502), .B2(new_n462), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n498), .B(G2104), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n494), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n505), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n491), .B2(new_n493), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT72), .A3(new_n504), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n518), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT74), .ZN(new_n521));
  OAI21_X1  g096(.A(G651), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT6), .B(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n523), .A3(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT73), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT73), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n530), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n518), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n523), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  INV_X1    g121(.A(new_n517), .ZN(new_n547));
  NOR2_X1   g122(.A1(KEYINPUT5), .A2(G543), .ZN(new_n548));
  AND2_X1   g123(.A1(KEYINPUT6), .A2(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n547), .A2(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n535), .A2(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n545), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n544), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n535), .A2(new_n557), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(new_n535), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n566), .A2(KEYINPUT76), .A3(G53), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n535), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n538), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n551), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n574), .A2(G651), .B1(G91), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n571), .B(new_n576), .C1(KEYINPUT9), .C2(new_n570), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n575), .A2(G87), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n535), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n581), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n566), .A2(G49), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n588), .A2(new_n582), .A3(KEYINPUT77), .A4(new_n584), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n516), .B2(new_n517), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n518), .A2(new_n523), .A3(G86), .ZN(new_n597));
  OAI211_X1 g172(.A(G48), .B(G543), .C1(new_n549), .C2(new_n550), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n544), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT78), .B(G85), .Z(new_n603));
  OAI22_X1  g178(.A1(new_n535), .A2(new_n602), .B1(new_n551), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n575), .A2(G92), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n538), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(G54), .B2(new_n566), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n607), .B1(new_n616), .B2(G868), .ZN(G321));
  XNOR2_X1  g192(.A(G321), .B(KEYINPUT80), .ZN(G284));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G297));
  XNOR2_X1  g196(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n615), .A2(G559), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n625), .A2(KEYINPUT82), .A3(new_n619), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT82), .B1(new_n625), .B2(new_n619), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n626), .B(new_n627), .C1(G868), .C2(new_n560), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g204(.A1(new_n478), .A2(new_n469), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n630), .B(new_n631), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n481), .A2(G123), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G135), .B2(new_n479), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n636), .A2(new_n637), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n655), .ZN(G401));
  INV_X1    g237(.A(KEYINPUT18), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2100), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(G2096), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n671), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n679), .B1(new_n681), .B2(new_n683), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n681), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n688), .C1(new_n678), .C2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(G303), .A2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G1971), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n697), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(G6), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n597), .A2(new_n598), .ZN(new_n705));
  OAI21_X1  g280(.A(G61), .B1(new_n547), .B2(new_n548), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n544), .B1(new_n706), .B2(new_n594), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n704), .B1(new_n708), .B2(new_n698), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n698), .A2(G23), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n583), .A2(new_n586), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n698), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  NAND4_X1  g291(.A1(new_n701), .A2(new_n703), .A3(new_n711), .A4(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n479), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n481), .A2(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n462), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT35), .B(G1991), .Z(new_n729));
  AND2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n698), .A2(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n605), .B2(new_n698), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1986), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n718), .A2(new_n719), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT36), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n718), .A2(new_n738), .A3(new_n719), .A4(new_n735), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT92), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT25), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(G127), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n478), .B2(new_n745), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n746), .A2(G2105), .B1(new_n479), .B2(G139), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G33), .B(new_n748), .S(G29), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2072), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n479), .A2(G141), .ZN(new_n752));
  INV_X1    g327(.A(G105), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(new_n469), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n481), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n720), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n720), .A2(G32), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n760), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n762), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n642), .A2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT30), .B(G28), .ZN(new_n767));
  OR2_X1    g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  NAND2_X1  g343(.A1(KEYINPUT31), .A2(G11), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n767), .A2(new_n720), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(G168), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G21), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT95), .B(G1966), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n764), .A2(new_n765), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G5), .A2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT96), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G301), .B2(new_n698), .ZN(new_n779));
  INV_X1    g354(.A(G1961), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n773), .B2(new_n774), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n720), .B1(new_n784), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G160), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2084), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n776), .A2(new_n782), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n720), .A2(G27), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G164), .B2(new_n720), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(new_n444), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n751), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n751), .A2(KEYINPUT97), .A3(new_n789), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n698), .A2(G20), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT23), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT100), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT99), .B(G1956), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G162), .A2(G29), .ZN(new_n803));
  OR2_X1    g378(.A1(G29), .A2(G35), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  INV_X1    g384(.A(G2090), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G4), .A2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT91), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n615), .B2(new_n698), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1348), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n720), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT28), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n479), .A2(G140), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n481), .A2(G128), .ZN(new_n819));
  OR2_X1    g394(.A1(G104), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(new_n720), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G2067), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n698), .A2(G19), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n560), .B2(new_n698), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1341), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n810), .B1(new_n808), .B2(new_n809), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n811), .A2(new_n815), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n802), .A2(new_n831), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n795), .A2(new_n796), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n740), .A2(new_n833), .ZN(G311));
  AND3_X1   g409(.A1(new_n833), .A2(new_n740), .A3(KEYINPUT101), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT101), .B1(new_n833), .B2(new_n740), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(G150));
  NAND2_X1  g412(.A1(new_n616), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n544), .ZN(new_n841));
  INV_X1    g416(.A(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI22_X1  g418(.A1(new_n535), .A2(new_n842), .B1(new_n551), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n560), .A2(new_n845), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n556), .A2(new_n559), .B1(new_n841), .B2(new_n844), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n839), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT102), .Z(new_n853));
  OAI21_X1  g428(.A(G860), .B1(new_n841), .B2(new_n844), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  NAND3_X1  g431(.A1(new_n743), .A2(KEYINPUT104), .A3(new_n747), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n759), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n506), .A2(KEYINPUT103), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n510), .A2(new_n860), .A3(new_n504), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n858), .B(new_n862), .Z(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n726), .B(KEYINPUT105), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n479), .A2(G142), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n462), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n865), .A2(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(new_n632), .ZN(new_n873));
  OR3_X1    g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n822), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n822), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n864), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n876), .A3(new_n863), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n642), .B(G160), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(G395));
  XNOR2_X1  g465(.A(new_n625), .B(new_n848), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n615), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n615), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  XOR2_X1   g471(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n891), .B(new_n899), .C1(KEYINPUT41), .C2(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n605), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n708), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(G166), .A2(new_n713), .ZN(new_n907));
  NOR2_X1   g482(.A1(G166), .A2(new_n713), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n905), .B1(new_n908), .B2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n896), .A2(new_n900), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n902), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n902), .B2(new_n915), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n845), .A2(G868), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n902), .A2(new_n915), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n912), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n619), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n919), .B2(new_n921), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(G331));
  NAND2_X1  g504(.A1(new_n848), .A2(G171), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n846), .A2(G301), .A3(new_n847), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(G286), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(G286), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n897), .B1(new_n892), .B2(new_n893), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n935), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n895), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n912), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n940), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n943), .B2(new_n913), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n912), .B1(new_n938), .B2(new_n940), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT109), .B1(new_n947), .B2(G37), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT43), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n940), .A2(KEYINPUT110), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n894), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n892), .A2(new_n893), .A3(new_n898), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n934), .A2(new_n935), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n940), .A2(KEYINPUT110), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n913), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND4_X1   g532(.A1(KEYINPUT43), .A2(new_n957), .A3(new_n885), .A4(new_n941), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n949), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n946), .B2(new_n948), .ZN(new_n962));
  AND4_X1   g537(.A1(new_n961), .A2(new_n957), .A3(new_n885), .A4(new_n941), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n862), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G125), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT3), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n467), .ZN(new_n972));
  NAND2_X1  g547(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n475), .B1(new_n974), .B2(new_n473), .ZN(new_n975));
  INV_X1    g550(.A(new_n474), .ZN(new_n976));
  OAI21_X1  g551(.A(G2105), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n470), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(G40), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n969), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n822), .B(G2067), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n759), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n729), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n726), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n980), .ZN(new_n989));
  NOR2_X1   g564(.A1(G290), .A2(G1986), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT111), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(G1986), .B2(G290), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT112), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n995));
  INV_X1    g570(.A(G1966), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n997), .B(new_n470), .C1(new_n476), .C2(G2105), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n510), .B2(new_n504), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n968), .A2(G1384), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n508), .B2(new_n511), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n995), .B(new_n996), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n979), .B1(new_n1005), .B2(new_n999), .ZN(new_n1006));
  INV_X1    g581(.A(G2084), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1384), .B1(new_n508), .B2(new_n511), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n506), .B2(new_n966), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n979), .ZN(new_n1012));
  AND4_X1   g587(.A1(KEYINPUT72), .A2(new_n494), .A3(new_n504), .A4(new_n505), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT72), .B1(new_n510), .B2(new_n504), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1001), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n995), .B1(new_n1016), .B2(new_n996), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G286), .A2(G8), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT123), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1021), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT51), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n996), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT118), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1009), .A3(new_n1004), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1023), .B1(new_n1028), .B2(G8), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1022), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n859), .A2(new_n861), .A3(new_n1001), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n859), .A2(KEYINPUT113), .A3(new_n861), .A4(new_n1001), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n966), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n979), .B1(new_n1036), .B2(new_n968), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1971), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1008), .A2(new_n1005), .ZN(new_n1039));
  INV_X1    g614(.A(new_n999), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n979), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1039), .A2(new_n1041), .A3(new_n810), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n529), .A2(G8), .A3(new_n531), .ZN(new_n1044));
  XOR2_X1   g619(.A(new_n1044), .B(KEYINPUT55), .Z(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(G305), .B2(G1981), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n707), .B1(new_n705), .B2(KEYINPUT116), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n597), .A2(new_n1050), .A3(new_n598), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1048), .B1(new_n1052), .B2(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  AOI211_X1 g629(.A(KEYINPUT117), .B(new_n1054), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n708), .B2(new_n1054), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1051), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1050), .B1(new_n597), .B2(new_n598), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n707), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(new_n1054), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1052), .A2(new_n1058), .A3(G1981), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT49), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(G160), .A2(G40), .A3(new_n506), .A4(new_n966), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(new_n1067), .A3(G8), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1066), .B2(G8), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1057), .A2(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n713), .A2(G1976), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT115), .B(G1976), .Z(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1071), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1070), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1005), .B1(new_n512), .B2(new_n966), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n998), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1078), .A2(new_n1079), .A3(G2090), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1045), .B(G8), .C1(new_n1038), .C2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1047), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1030), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1035), .A2(new_n1037), .A3(new_n444), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1006), .B(KEYINPUT120), .C1(new_n1008), .C2(new_n1005), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n780), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1012), .A2(new_n1015), .A3(new_n444), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1012), .A2(new_n1015), .A3(KEYINPUT124), .A4(new_n444), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1086), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n979), .A2(KEYINPUT125), .ZN(new_n1099));
  NOR4_X1   g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n1085), .A4(G2078), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(new_n1035), .A3(new_n969), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1086), .A2(new_n1090), .A3(new_n1101), .A4(G301), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1086), .A2(new_n1090), .A3(new_n1101), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G171), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(KEYINPUT54), .C1(G171), .C2(new_n1096), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1083), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  XOR2_X1   g684(.A(G299), .B(KEYINPUT57), .Z(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1035), .A2(new_n1037), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1113));
  INV_X1    g688(.A(G1956), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1115), .A3(new_n1110), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT61), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1066), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT58), .B(G1341), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1035), .A2(new_n1037), .A3(new_n982), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(KEYINPUT121), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(KEYINPUT121), .B2(new_n1125), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n560), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1088), .A2(new_n1131), .A3(new_n1089), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1066), .A2(G2067), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT119), .Z(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1134), .A3(KEYINPUT60), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT60), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(new_n615), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1132), .A2(new_n1134), .A3(KEYINPUT60), .A4(new_n616), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1129), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1127), .A2(new_n560), .A3(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1121), .A2(new_n1130), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n615), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1116), .B1(new_n1143), .B2(new_n1118), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1109), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1030), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT51), .A3(new_n1024), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1150), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1022), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1030), .A2(new_n1147), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1082), .A2(new_n1097), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NOR4_X1   g729(.A1(new_n1057), .A2(new_n1065), .A3(G1976), .A4(G288), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G305), .A2(G1981), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1155), .A2(new_n1156), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1077), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1081), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT63), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1028), .A2(G8), .A3(G168), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1082), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1160), .ZN(new_n1163));
  OAI21_X1  g738(.A(G8), .B1(new_n1038), .B2(new_n1080), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1046), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1163), .A2(new_n1081), .A3(new_n1077), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1159), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n994), .B1(new_n1145), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n759), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n980), .B1(new_n1170), .B2(new_n981), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n980), .A2(new_n982), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1172), .A2(KEYINPUT46), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(KEYINPUT46), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT47), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n980), .A2(new_n991), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT48), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n988), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n822), .A2(G2067), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n727), .A2(new_n985), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n984), .B2(new_n1183), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1180), .A2(new_n1181), .B1(new_n989), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1176), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1169), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n1189));
  AND3_X1   g763(.A1(new_n675), .A2(KEYINPUT127), .A3(new_n460), .ZN(new_n1190));
  AOI21_X1  g764(.A(KEYINPUT127), .B1(new_n675), .B2(new_n460), .ZN(new_n1191));
  NOR4_X1   g765(.A1(G229), .A2(new_n1190), .A3(new_n1191), .A4(G401), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n886), .B2(new_n887), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1189), .A2(new_n1193), .ZN(G308));
  OAI221_X1 g768(.A(new_n1192), .B1(new_n887), .B2(new_n886), .C1(new_n962), .C2(new_n963), .ZN(G225));
endmodule


