//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n254, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n261, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(KEYINPUT66), .A2(G68), .ZN(new_n214));
  NOR2_X1   g0014(.A1(KEYINPUT66), .A2(G68), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n218), .B(new_n222), .C1(new_n227), .C2(KEYINPUT68), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n213), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT69), .ZN(new_n233));
  INV_X1    g0033(.A(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n213), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n236), .B(G250), .C1(G257), .C2(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT0), .ZN(new_n238));
  NAND2_X1  g0038(.A1(G1), .A2(G13), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G20), .ZN(new_n241));
  INV_X1    g0041(.A(new_n203), .ZN(new_n242));
  OR2_X1    g0042(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n243), .A2(G50), .A3(new_n244), .ZN(new_n245));
  OAI221_X1 g0045(.A(new_n238), .B1(new_n241), .B2(new_n245), .C1(new_n230), .C2(new_n231), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n233), .A2(new_n246), .ZN(G361));
  XNOR2_X1  g0047(.A(G238), .B(G244), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G232), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT2), .B(G226), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G264), .B(G270), .Z(new_n252));
  XNOR2_X1  g0052(.A(G250), .B(G257), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G358));
  XNOR2_X1  g0055(.A(G50), .B(G68), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G58), .B(G77), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n256), .B(new_n257), .Z(new_n258));
  XNOR2_X1  g0058(.A(G87), .B(G97), .ZN(new_n259));
  XNOR2_X1  g0059(.A(G107), .B(G116), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n258), .B(new_n261), .Z(G351));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n239), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT71), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n263), .A2(new_n266), .A3(new_n239), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n234), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n211), .B2(G20), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n272), .A2(new_n274), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(G58), .B1(new_n214), .B2(new_n215), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT74), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(KEYINPUT74), .B(G58), .C1(new_n214), .C2(new_n215), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n203), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G159), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n212), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT7), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n287), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n216), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n282), .A2(new_n284), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT16), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n264), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n281), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n293), .B2(G68), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n276), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G41), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n240), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n239), .B1(G33), .B2(G41), .ZN(new_n311));
  INV_X1    g0111(.A(G41), .ZN(new_n312));
  INV_X1    g0112(.A(G45), .ZN(new_n313));
  AOI21_X1  g0113(.A(G1), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G232), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  INV_X1    g0118(.A(new_n311), .ZN(new_n319));
  INV_X1    g0119(.A(G226), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G1698), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n321), .B1(G223), .B2(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G87), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n317), .A2(new_n318), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n307), .B(KEYINPUT70), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n306), .B1(new_n315), .B2(G232), .ZN(new_n330));
  INV_X1    g0130(.A(new_n326), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT18), .B1(new_n303), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n301), .A2(new_n282), .A3(new_n284), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n264), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT16), .B1(new_n300), .B2(new_n295), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n275), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  INV_X1    g0139(.A(new_n333), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G200), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n317), .B2(new_n326), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n330), .A2(new_n331), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n275), .B(new_n346), .C1(new_n336), .C2(new_n337), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT17), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n303), .A2(KEYINPUT17), .A3(new_n346), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n334), .A2(new_n341), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n310), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G226), .B2(new_n315), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n287), .A2(new_n288), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(new_n220), .B2(new_n355), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n322), .A2(new_n323), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(G222), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n354), .B1(new_n319), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n211), .A2(G20), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n272), .A2(G50), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n283), .A2(G150), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n212), .A2(G33), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n273), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G50), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n212), .B1(new_n242), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n268), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n271), .A2(new_n368), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n364), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n362), .A2(G200), .B1(new_n373), .B2(KEYINPUT9), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(KEYINPUT9), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n344), .C2(new_n362), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT10), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n362), .B2(new_n328), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(G179), .B2(new_n362), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n283), .A2(G50), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n381), .B1(new_n220), .B2(new_n366), .C1(new_n294), .C2(new_n212), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n268), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT11), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT12), .B1(new_n294), .B2(new_n270), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  OR3_X1    g0189(.A1(new_n270), .A2(KEYINPUT12), .A3(G68), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n271), .A2(new_n264), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G68), .A3(new_n363), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n382), .A2(KEYINPUT11), .A3(new_n268), .ZN(new_n394));
  AND4_X1   g0194(.A1(new_n385), .A2(new_n391), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n329), .A2(new_n306), .B1(new_n315), .B2(G238), .ZN(new_n396));
  INV_X1    g0196(.A(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n320), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n355), .B(new_n398), .C1(G232), .C2(new_n397), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G97), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n319), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI211_X1 g0203(.A(KEYINPUT72), .B(new_n319), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n396), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n396), .C1(new_n403), .C2(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n395), .B1(new_n409), .B2(new_n344), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n342), .B1(new_n406), .B2(new_n408), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(G179), .A3(new_n408), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n409), .A2(new_n416), .A3(G169), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n395), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n412), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n360), .A2(G232), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n206), .B2(new_n355), .C1(new_n217), .C2(new_n356), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n311), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n353), .B1(G244), .B2(new_n315), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n392), .A2(G77), .A3(new_n363), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(G77), .B2(new_n270), .ZN(new_n428));
  INV_X1    g0228(.A(new_n273), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n429), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(new_n366), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n299), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n426), .B(new_n434), .C1(new_n344), .C2(new_n425), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n425), .A2(new_n328), .ZN(new_n437));
  INV_X1    g0237(.A(new_n434), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n423), .A2(new_n318), .A3(new_n424), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n352), .A2(new_n380), .A3(new_n420), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n271), .A2(new_n206), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT25), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n211), .A2(G33), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n265), .A2(new_n270), .A3(new_n267), .A4(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n206), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n355), .A2(new_n212), .A3(G87), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT22), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT23), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n212), .B2(G107), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n454), .A2(new_n455), .B1(new_n457), .B2(new_n212), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT24), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n452), .A2(new_n461), .A3(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n450), .B1(new_n463), .B2(new_n264), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT81), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n355), .A2(G257), .A3(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G294), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n355), .A2(new_n397), .ZN(new_n468));
  INV_X1    g0268(.A(G250), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT80), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n311), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n313), .A2(G1), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n319), .A3(G264), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n306), .A2(new_n474), .A3(new_n473), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n471), .B1(new_n470), .B2(new_n311), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n465), .B(G169), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n477), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(KEYINPUT82), .B2(new_n476), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n311), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n476), .A2(KEYINPUT82), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(G179), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n480), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n472), .A3(new_n478), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G169), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT81), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n464), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n342), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n489), .B2(G190), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n464), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n355), .A2(G250), .A3(G1698), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n355), .A2(G244), .A3(new_n397), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT4), .B1(new_n360), .B2(G244), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n311), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n311), .B1(new_n474), .B2(new_n473), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n482), .B1(G257), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n270), .A2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n447), .B2(new_n205), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n293), .A2(G107), .ZN(new_n512));
  OR2_X1    g0312(.A1(KEYINPUT76), .A2(G97), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT76), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(G107), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G97), .A2(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n207), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G20), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n283), .A2(G77), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT75), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n512), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n511), .B1(new_n527), .B2(new_n264), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n508), .B(new_n528), .C1(new_n344), .C2(new_n507), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n515), .A2(new_n517), .B1(new_n520), .B2(new_n516), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n530), .B2(new_n212), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n206), .B1(new_n291), .B2(new_n292), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n264), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n511), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n504), .A2(new_n506), .A3(new_n318), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n504), .A2(new_n506), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(G169), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n529), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT77), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n529), .A2(new_n541), .A3(new_n538), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n355), .A2(G264), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n355), .A2(G257), .A3(new_n397), .ZN(new_n545));
  INV_X1    g0345(.A(G303), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n355), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n311), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(KEYINPUT79), .A3(new_n311), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n498), .A2(new_n212), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n515), .B2(new_n286), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n264), .A2(new_n557), .ZN(new_n558));
  OR3_X1    g0358(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n555), .B1(new_n554), .B2(new_n558), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n211), .B2(G33), .ZN(new_n562));
  INV_X1    g0362(.A(new_n557), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n392), .A2(new_n562), .B1(new_n269), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n505), .A2(G270), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n477), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n552), .A2(new_n565), .A3(G179), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n551), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT79), .B1(new_n547), .B2(new_n311), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n328), .B1(new_n561), .B2(new_n564), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n569), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n552), .A2(G190), .A3(new_n568), .ZN(new_n578));
  INV_X1    g0378(.A(new_n565), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n567), .B1(new_n550), .B2(new_n551), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n579), .C1(new_n342), .C2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n355), .A2(new_n212), .A3(G68), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n366), .B1(new_n513), .B2(new_n514), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(KEYINPUT19), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n586), .A2(new_n212), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n513), .A2(new_n514), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G87), .A2(G107), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n264), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n271), .A2(new_n431), .ZN(new_n592));
  INV_X1    g0392(.A(G87), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n447), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n355), .A2(G244), .A3(G1698), .ZN(new_n596));
  OAI211_X1 g0396(.A(G238), .B(new_n397), .C1(new_n322), .C2(new_n323), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n456), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n311), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n311), .A2(new_n469), .A3(new_n474), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n306), .B2(new_n474), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n601), .A3(G190), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n599), .A2(new_n601), .A3(KEYINPUT78), .A4(G190), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n601), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n595), .A2(new_n604), .A3(new_n605), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n328), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n447), .A2(new_n431), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n591), .A2(new_n592), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n599), .A2(new_n601), .A3(new_n318), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n577), .A2(new_n582), .A3(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n443), .A2(new_n497), .A3(new_n543), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT83), .ZN(G372));
  OAI21_X1  g0417(.A(KEYINPUT26), .B1(new_n614), .B2(new_n538), .ZN(new_n618));
  INV_X1    g0418(.A(new_n536), .ZN(new_n619));
  AOI21_X1  g0419(.A(G169), .B1(new_n504), .B2(new_n506), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n619), .A2(new_n528), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT19), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n588), .B2(new_n366), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n515), .A2(G87), .A3(G107), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n583), .C1(new_n625), .C2(new_n587), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n264), .B1(new_n271), .B2(new_n431), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n607), .A2(new_n627), .A3(new_n602), .A4(new_n594), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n621), .A2(new_n622), .A3(new_n613), .A4(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n618), .A2(new_n613), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n539), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n613), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n464), .B2(new_n495), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n631), .B(new_n633), .C1(new_n492), .C2(new_n577), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n443), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n412), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n349), .A3(new_n350), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n417), .A2(new_n415), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n416), .B1(new_n409), .B2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n419), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n440), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n334), .A2(new_n341), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n377), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n379), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n636), .A2(new_n645), .ZN(G369));
  INV_X1    g0446(.A(new_n577), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n269), .A2(new_n212), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n647), .B(new_n581), .C1(new_n579), .C2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n577), .A2(new_n565), .A3(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n497), .B1(new_n464), .B2(new_n654), .ZN(new_n660));
  INV_X1    g0460(.A(new_n492), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n654), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n647), .A2(new_n653), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n497), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n492), .A2(new_n654), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(G399));
  NAND2_X1  g0469(.A1(new_n625), .A2(new_n556), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n235), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G1), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n671), .A2(new_n674), .B1(new_n245), .B2(new_n673), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n653), .B1(new_n630), .B2(new_n634), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(KEYINPUT29), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n621), .A2(new_n622), .A3(new_n613), .A4(new_n608), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT26), .B1(new_n632), .B2(new_n538), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n613), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT86), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT86), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n680), .A2(new_n681), .A3(new_n684), .A4(new_n613), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n634), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n654), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n615), .A2(new_n497), .A3(new_n543), .A4(new_n654), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  INV_X1    g0491(.A(new_n606), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n537), .A2(new_n552), .A3(new_n566), .A4(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n691), .B1(new_n693), .B2(new_n486), .ZN(new_n694));
  INV_X1    g0494(.A(new_n566), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n695), .B(new_n606), .C1(new_n550), .C2(new_n551), .ZN(new_n696));
  INV_X1    g0496(.A(new_n486), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(KEYINPUT30), .A3(new_n697), .A4(new_n537), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n692), .A2(G179), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n572), .A3(new_n493), .A4(new_n507), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n694), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n653), .ZN(new_n702));
  XNOR2_X1  g0502(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n690), .B(new_n705), .C1(KEYINPUT31), .C2(new_n702), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n679), .B(new_n689), .C1(G330), .C2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n676), .B1(new_n707), .B2(G1), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT87), .ZN(G364));
  NOR2_X1   g0509(.A1(new_n234), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n211), .B1(new_n710), .B2(G45), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n673), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n659), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G330), .B2(new_n657), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n239), .B1(G20), .B2(new_n328), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n212), .A2(new_n342), .A3(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G190), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n212), .A2(new_n318), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(G190), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(G326), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n719), .A2(new_n546), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(G200), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G190), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(KEYINPUT33), .A2(G317), .ZN(new_n727));
  NAND2_X1  g0527(.A1(KEYINPUT33), .A2(G317), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n212), .B1(new_n730), .B2(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n723), .B(new_n729), .C1(G294), .C2(new_n732), .ZN(new_n733));
  NOR4_X1   g0533(.A1(new_n212), .A2(new_n318), .A3(G190), .A4(G200), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT89), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G311), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n730), .A2(G20), .A3(new_n344), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT90), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G329), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n342), .A2(G20), .A3(G179), .A4(G190), .ZN(new_n746));
  INV_X1    g0546(.A(G322), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n359), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n718), .A2(new_n344), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(G283), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n733), .A2(new_n739), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n731), .A2(new_n205), .ZN(new_n753));
  INV_X1    g0553(.A(new_n740), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G159), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n755), .A2(KEYINPUT32), .B1(new_n719), .B2(new_n593), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n753), .B(new_n756), .C1(G68), .C2(new_n725), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n738), .A2(G77), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n749), .A2(new_n206), .ZN(new_n759));
  INV_X1    g0559(.A(new_n746), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n359), .B(new_n759), .C1(G58), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n721), .ZN(new_n762));
  AOI22_X1  g0562(.A1(KEYINPUT32), .A2(new_n755), .B1(new_n762), .B2(G50), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n757), .A2(new_n758), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n717), .B1(new_n752), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n236), .A2(new_n355), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n209), .A2(new_n766), .B1(G116), .B2(new_n236), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n235), .A2(new_n355), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT88), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n245), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n313), .B2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n258), .A2(new_n313), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n767), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n716), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n713), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n765), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n777), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n657), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n715), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  NAND2_X1  g0585(.A1(new_n440), .A2(KEYINPUT93), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT93), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n437), .A2(new_n787), .A3(new_n438), .A4(new_n439), .ZN(new_n788));
  AND3_X1   g0588(.A1(new_n786), .A2(new_n435), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n677), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n438), .A2(new_n653), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n435), .A3(new_n791), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n441), .A2(new_n653), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n790), .B1(new_n677), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n706), .A2(G330), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT94), .Z(new_n799));
  AOI21_X1  g0599(.A(new_n713), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n717), .A2(new_n776), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n713), .B1(G77), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n749), .A2(new_n593), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n726), .A2(new_n805), .B1(new_n721), .B2(new_n546), .ZN(new_n806));
  INV_X1    g0606(.A(new_n719), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n806), .C1(G107), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n744), .A2(G311), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n738), .A2(G116), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n355), .B(new_n753), .C1(G294), .C2(new_n760), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n762), .A2(G137), .B1(G143), .B2(new_n760), .ZN(new_n813));
  INV_X1    g0613(.A(G150), .ZN(new_n814));
  INV_X1    g0614(.A(new_n738), .ZN(new_n815));
  INV_X1    g0615(.A(G159), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n813), .B1(new_n814), .B2(new_n726), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT34), .Z(new_n818));
  AOI22_X1  g0618(.A1(new_n807), .A2(G50), .B1(new_n732), .B2(G58), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n359), .B1(new_n750), .B2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n743), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT91), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n812), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT92), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n717), .B1(new_n824), .B2(KEYINPUT92), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n803), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n776), .B2(new_n795), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n801), .A2(new_n828), .ZN(G384));
  AOI211_X1 g0629(.A(new_n556), .B(new_n241), .C1(new_n522), .C2(KEYINPUT35), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(KEYINPUT35), .B2(new_n522), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT36), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n771), .A2(G77), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n279), .A2(new_n280), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(G50), .B2(new_n202), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n835), .A2(G1), .A3(new_n234), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT95), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n293), .A2(G68), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n282), .A2(new_n284), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n297), .ZN(new_n841));
  INV_X1    g0641(.A(new_n268), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n300), .B2(new_n301), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n276), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n347), .B(KEYINPUT96), .C1(new_n333), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n335), .A2(new_n268), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT16), .B1(new_n300), .B2(new_n839), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n275), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n651), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n340), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT96), .B1(new_n852), .B2(new_n347), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT97), .B1(new_n303), .B2(new_n651), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT97), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n338), .A2(new_n856), .A3(new_n849), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n347), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n298), .A2(new_n302), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n333), .B1(new_n860), .B2(new_n275), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n850), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n854), .A2(new_n864), .B1(new_n351), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n419), .A2(new_n653), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n641), .A2(new_n637), .A3(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n419), .B(new_n653), .C1(new_n418), .C2(new_n412), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n653), .B1(new_n786), .B2(new_n788), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n677), .B2(new_n789), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n869), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n643), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n849), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT99), .ZN(new_n880));
  INV_X1    g0680(.A(new_n858), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n351), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n858), .A2(new_n862), .A3(new_n863), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n863), .B1(new_n858), .B2(new_n862), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(KEYINPUT98), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT98), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n868), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n880), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT98), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n858), .A2(new_n862), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n896), .A2(new_n864), .B1(new_n351), .B2(new_n881), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n894), .B1(new_n897), .B2(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n885), .A2(KEYINPUT98), .A3(new_n886), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(KEYINPUT99), .A3(new_n890), .A4(new_n868), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n892), .A2(new_n893), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n418), .A2(new_n419), .A3(new_n654), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n879), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n443), .B1(new_n689), .B2(new_n679), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n645), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n905), .B(new_n907), .Z(new_n908));
  INV_X1    g0708(.A(G330), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n794), .B1(new_n871), .B2(new_n872), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n704), .B1(new_n701), .B2(new_n653), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n690), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT40), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n868), .B1(new_n887), .B2(new_n888), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT100), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT100), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n900), .A2(new_n919), .A3(new_n868), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n869), .A2(new_n915), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n443), .A2(new_n914), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n908), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n211), .B2(new_n710), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n908), .A2(new_n927), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n838), .B1(new_n929), .B2(new_n930), .ZN(G367));
  OAI21_X1  g0731(.A(new_n631), .B1(new_n528), .B2(new_n654), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n621), .A2(new_n653), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT101), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n492), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n653), .B1(new_n937), .B2(new_n538), .ZN(new_n938));
  INV_X1    g0738(.A(new_n934), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n665), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n595), .A2(new_n654), .ZN(new_n943));
  MUX2_X1   g0743(.A(new_n632), .B(new_n613), .S(new_n943), .Z(new_n944));
  OAI22_X1  g0744(.A1(new_n938), .A2(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n942), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n663), .A2(new_n935), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n672), .B(KEYINPUT41), .Z(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n668), .B2(new_n934), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT103), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n939), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT102), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n955), .A2(new_n956), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n667), .A2(new_n939), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n663), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n665), .B1(new_n662), .B2(new_n664), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n659), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n707), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n961), .A2(new_n663), .A3(new_n963), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n965), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n951), .B1(new_n971), .B2(new_n707), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n711), .B(KEYINPUT104), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n949), .B(new_n950), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(G137), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n355), .B1(new_n746), .B2(new_n814), .C1(new_n740), .C2(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n726), .A2(new_n816), .B1(new_n220), .B2(new_n749), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G50), .C2(new_n738), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n807), .A2(G58), .B1(new_n762), .B2(G143), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n202), .C2(new_n731), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n807), .A2(G116), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n359), .B1(new_n746), .B2(new_n546), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G317), .B2(new_n754), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n805), .C2(new_n815), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n762), .A2(G311), .B1(new_n732), .B2(G107), .ZN(new_n986));
  INV_X1    g0786(.A(G294), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n986), .B1(new_n588), .B2(new_n749), .C1(new_n987), .C2(new_n726), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n980), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n716), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n944), .A2(new_n777), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n778), .B1(new_n236), .B2(new_n431), .C1(new_n770), .C2(new_n254), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n991), .A2(new_n713), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n974), .A2(new_n994), .ZN(G387));
  OAI21_X1  g0795(.A(new_n769), .B1(new_n251), .B2(new_n313), .ZN(new_n996));
  INV_X1    g0796(.A(new_n671), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n997), .B2(new_n766), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n313), .B1(new_n202), .B2(new_n220), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n429), .A2(new_n368), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n997), .B(new_n1001), .C1(KEYINPUT50), .C2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n998), .A2(new_n1002), .B1(new_n206), .B2(new_n235), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n713), .B1(new_n1003), .B2(new_n779), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n355), .B1(new_n740), .B2(new_n814), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n726), .A2(new_n273), .B1(new_n816), .B2(new_n721), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G50), .C2(new_n760), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n731), .A2(new_n431), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n719), .A2(new_n220), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G97), .C2(new_n750), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1007), .B(new_n1010), .C1(new_n202), .C2(new_n815), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n355), .B1(new_n754), .B2(G326), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n807), .A2(G294), .B1(new_n732), .B2(G283), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n725), .A2(G311), .B1(G317), .B2(new_n760), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n747), .B2(new_n721), .C1(new_n815), .C2(new_n546), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT105), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1013), .B1(new_n1017), .B2(KEYINPUT48), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT48), .B2(new_n1017), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT106), .Z(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1012), .B1(new_n556), .B2(new_n749), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1011), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1004), .B1(new_n1024), .B2(new_n716), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n662), .A2(new_n782), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n1026), .B1(new_n967), .B2(new_n973), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n969), .A2(new_n673), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n707), .B2(new_n967), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(G393));
  INV_X1    g0830(.A(new_n970), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n968), .B1(new_n1031), .B2(new_n964), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1032), .A2(new_n971), .A3(new_n672), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n965), .A2(new_n970), .A3(new_n973), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n726), .A2(new_n546), .B1(new_n731), .B2(new_n556), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G283), .B2(new_n807), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n355), .B(new_n759), .C1(G322), .C2(new_n754), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n987), .C2(new_n815), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n762), .A2(G317), .B1(G311), .B2(new_n760), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n721), .A2(new_n814), .B1(new_n816), .B2(new_n746), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT51), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n726), .A2(new_n368), .B1(new_n731), .B2(new_n220), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n294), .B2(new_n807), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n359), .B(new_n804), .C1(G143), .C2(new_n754), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n738), .A2(new_n429), .ZN(new_n1048));
  AND4_X1   g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n716), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n769), .A2(new_n261), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n779), .B1(new_n235), .B2(new_n515), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n712), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT107), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1050), .B(new_n1054), .C1(new_n936), .C2(new_n782), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1033), .A2(new_n1034), .A3(new_n1055), .ZN(G390));
  AOI21_X1  g0856(.A(new_n909), .B1(new_n913), .B2(new_n690), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n443), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n906), .A2(new_n645), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n686), .A2(new_n654), .A3(new_n789), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n874), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT109), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(KEYINPUT109), .A3(new_n1061), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n706), .A2(G330), .A3(new_n795), .A4(new_n873), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n909), .B(new_n794), .C1(new_n913), .C2(new_n690), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n873), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n873), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n797), .B2(new_n794), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1057), .A2(new_n910), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n875), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1059), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1064), .A2(new_n873), .A3(new_n1065), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n919), .B1(new_n900), .B2(new_n868), .ZN(new_n1077));
  AOI221_X4 g0877(.A(new_n886), .B1(new_n351), .B2(new_n865), .C1(new_n854), .C2(new_n864), .ZN(new_n1078));
  AOI211_X1 g0878(.A(KEYINPUT100), .B(new_n1078), .C1(new_n898), .C2(new_n899), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1076), .B(new_n903), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n903), .B1(new_n875), .B2(new_n1071), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n892), .A2(new_n901), .A3(new_n1081), .A4(new_n893), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1080), .A2(new_n1082), .A3(new_n1067), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1073), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1075), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1073), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n1082), .A3(new_n1067), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n906), .A2(new_n645), .A3(new_n1058), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1074), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n1067), .C1(new_n873), .C2(new_n1068), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1085), .A2(new_n1095), .A3(new_n672), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n355), .B1(new_n760), .B2(G116), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1097), .B1(new_n593), .B2(new_n719), .C1(new_n743), .C2(new_n987), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n750), .A2(G68), .B1(G77), .B2(new_n732), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n206), .B2(new_n726), .C1(new_n805), .C2(new_n721), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n515), .C2(new_n738), .ZN(new_n1101));
  INV_X1    g0901(.A(G125), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n355), .B1(new_n368), .B2(new_n749), .C1(new_n743), .C2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT110), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n815), .A2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n762), .A2(G128), .B1(G132), .B2(new_n760), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n816), .B2(new_n731), .C1(new_n975), .C2(new_n726), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT53), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n807), .B2(G150), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n719), .A2(KEYINPUT53), .A3(new_n814), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1101), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n713), .B1(new_n429), .B2(new_n802), .C1(new_n1113), .C2(new_n717), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n902), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n775), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n973), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1096), .A2(new_n1118), .ZN(G378));
  NAND2_X1  g0919(.A1(new_n910), .A2(new_n914), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n867), .B2(new_n868), .ZN(new_n1121));
  OAI21_X1  g0921(.A(G330), .B1(new_n1121), .B2(KEYINPUT40), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT114), .B1(new_n921), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1120), .A2(new_n922), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n909), .B1(new_n923), .B2(new_n922), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n372), .A2(new_n849), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT112), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n380), .B(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1123), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1125), .A2(new_n1133), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n905), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1135), .A2(new_n905), .A3(new_n1136), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n973), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n713), .B1(G50), .B2(new_n802), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n726), .A2(new_n821), .B1(new_n721), .B2(new_n1102), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G150), .B2(new_n732), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1105), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n807), .A2(new_n1145), .B1(G128), .B2(new_n760), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n975), .C2(new_n815), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n750), .A2(G159), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n749), .A2(new_n201), .B1(new_n721), .B2(new_n556), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1009), .B(new_n1153), .C1(G97), .C2(new_n725), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n355), .A2(G41), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n202), .B2(new_n731), .C1(new_n206), .C2(new_n746), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G283), .B2(new_n744), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1154), .B(new_n1157), .C1(new_n431), .C2(new_n815), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT58), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G50), .B(new_n1155), .C1(new_n286), .C2(new_n312), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT111), .Z(new_n1163));
  NAND4_X1  g0963(.A1(new_n1152), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1142), .B1(new_n1164), .B2(new_n716), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n1134), .B2(new_n776), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT113), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n1141), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT115), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1083), .A2(new_n1084), .A3(new_n1075), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n1090), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1095), .A2(KEYINPUT115), .A3(new_n1059), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1135), .A2(new_n905), .A3(new_n1136), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n905), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n672), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1169), .B1(new_n1180), .B2(new_n1182), .ZN(G375));
  OAI21_X1  g0983(.A(new_n713), .B1(G68), .B2(new_n802), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n726), .A2(new_n556), .B1(new_n721), .B2(new_n987), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1008), .B(new_n1185), .C1(G97), .C2(new_n807), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n744), .A2(G303), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n359), .B1(new_n746), .B2(new_n805), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n750), .B2(G77), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n738), .A2(G107), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n726), .A2(new_n1105), .B1(new_n368), .B2(new_n731), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n719), .A2(new_n816), .B1(new_n721), .B2(new_n821), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n738), .A2(G150), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n744), .A2(G128), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n355), .B1(new_n746), .B2(new_n975), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n750), .B2(G58), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT116), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n717), .B1(new_n1200), .B2(KEYINPUT116), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1184), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n873), .B2(new_n776), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n973), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1094), .A2(new_n951), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1090), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(G381));
  XOR2_X1   g1011(.A(G375), .B(KEYINPUT118), .Z(new_n1212));
  OR4_X1    g1012(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(G378), .B(KEYINPUT117), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(new_n1213), .A2(G387), .A3(new_n1214), .A4(G381), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(G407));
  AND2_X1   g1016(.A1(new_n1096), .A2(new_n1118), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT117), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n652), .A2(G213), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1212), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(G213), .A3(G407), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT119), .ZN(G409));
  NAND3_X1  g1023(.A1(new_n1205), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(new_n672), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1209), .B1(new_n1226), .B2(new_n1094), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1207), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G384), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(G384), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1095), .A2(KEYINPUT115), .A3(new_n1059), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT115), .B1(new_n1095), .B2(new_n1059), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1181), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1177), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n673), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1217), .B(new_n1168), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1141), .A2(new_n1166), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1175), .A2(new_n1176), .A3(new_n951), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1174), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(KEYINPUT120), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT120), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1174), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1214), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1219), .B(new_n1232), .C1(new_n1238), .C2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT121), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT63), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1247), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(G393), .B(new_n784), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n974), .A2(new_n994), .A3(G390), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G390), .B1(new_n974), .B2(new_n994), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1256), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1257), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1207), .ZN(new_n1265));
  INV_X1    g1065(.A(G2897), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1219), .A2(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1265), .A2(new_n1229), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1267), .B1(new_n1265), .B2(new_n1229), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1262), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1230), .A2(new_n1231), .B1(new_n1266), .B2(new_n1219), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1229), .A3(new_n1267), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(KEYINPUT122), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1219), .B1(new_n1238), .B2(new_n1245), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1261), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n951), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1139), .A2(new_n1279), .A3(new_n1140), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT120), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1239), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1244), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1218), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G378), .B(new_n1169), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1232), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n1248), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n1277), .A2(new_n1286), .A3(new_n1219), .A4(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1220), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1277), .B1(new_n1290), .B2(new_n1288), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1276), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT124), .B1(new_n1251), .B2(new_n1292), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1220), .B(new_n1287), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT121), .B1(new_n1294), .B2(KEYINPUT63), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT124), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1288), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT123), .B1(new_n1275), .B2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1290), .A2(new_n1277), .A3(new_n1288), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1297), .A2(new_n1298), .A3(new_n1302), .A4(new_n1276), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1293), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT125), .B1(new_n1294), .B2(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1294), .A2(new_n1306), .A3(KEYINPUT62), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT126), .B1(new_n1246), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT125), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1246), .A2(new_n1310), .A3(new_n1308), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1305), .A2(new_n1307), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1304), .A2(new_n1317), .ZN(G405));
  AOI21_X1  g1118(.A(new_n1238), .B1(G375), .B2(new_n1218), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT127), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1232), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1323), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1287), .A3(new_n1321), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1316), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1327), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


