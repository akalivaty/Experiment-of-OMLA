//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n447, new_n451, new_n452,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n451));
  AND2_X1   g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(G223));
  NAND2_X1  g028(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NOR4_X1   g032(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(new_n457), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(G2106), .B2(new_n464), .ZN(G319));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(G137), .A3(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n472), .A2(KEYINPUT69), .A3(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n472), .B2(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n469), .B1(new_n466), .B2(new_n467), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n476), .B2(new_n477), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n477), .C2(new_n476), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT70), .B1(new_n469), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(G126), .A2(new_n484), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n496), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .A3(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n511), .A2(new_n510), .B1(new_n522), .B2(new_n523), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(G651), .A2(new_n526), .B1(new_n528), .B2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n520), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  XOR2_X1   g106(.A(KEYINPUT73), .B(G89), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n518), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n539), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(G168));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n524), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n546), .B2(KEYINPUT74), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(KEYINPUT74), .B2(new_n546), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT75), .B(G90), .Z(new_n549));
  AOI22_X1  g124(.A1(new_n528), .A2(new_n549), .B1(new_n518), .B2(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n513), .A2(new_n553), .B1(new_n554), .B2(new_n527), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n539), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n513), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n518), .A2(new_n566), .A3(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n524), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(G651), .A2(new_n571), .B1(new_n528), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  XNOR2_X1  g148(.A(new_n541), .B(KEYINPUT76), .ZN(G286));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n513), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n518), .A2(KEYINPUT77), .A3(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n539), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n528), .B2(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n518), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n527), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n537), .B2(new_n538), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n512), .A2(new_n590), .A3(G86), .A4(new_n539), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n583), .A2(new_n585), .A3(new_n589), .A4(new_n591), .ZN(G305));
  XNOR2_X1  g167(.A(KEYINPUT79), .B(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n513), .A2(new_n593), .B1(new_n594), .B2(new_n527), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n539), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n528), .A2(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n513), .B2(KEYINPUT80), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n524), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n604), .A2(new_n606), .B1(G651), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G321));
  NOR2_X1   g188(.A1(G299), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n541), .B(KEYINPUT76), .Z(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  AOI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n468), .A2(new_n472), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT81), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n482), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n484), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n469), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2096), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n626), .B2(new_n627), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT83), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n644), .A2(new_n645), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n644), .A2(new_n645), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(G14), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n651), .A2(new_n656), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n661), .B2(new_n652), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  NOR3_X1   g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT17), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n667), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n673), .A2(new_n674), .A3(new_n666), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n666), .B2(new_n668), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n666), .B2(new_n673), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n670), .B(new_n675), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n627), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT87), .B(G2096), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n691), .B(new_n690), .S(new_n694), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n696));
  OR3_X1    g271(.A1(new_n687), .A2(new_n688), .A3(KEYINPUT89), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n695), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT91), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G303), .B2(G16), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G1971), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(G23), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n579), .A2(new_n581), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n710), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G6), .B(G305), .S(G16), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n714), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n482), .A2(G131), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G107), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n484), .A2(G119), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G29), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G25), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n710), .A2(G24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n598), .B2(new_n710), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1986), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n739), .B2(new_n740), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n726), .A2(new_n727), .A3(new_n741), .A4(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT36), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n558), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G19), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT98), .B(G1341), .Z(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G26), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT28), .Z(new_n754));
  AOI22_X1  g329(.A1(G128), .A2(new_n484), .B1(new_n482), .B2(G140), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n756), .A2(G104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(G104), .ZN(new_n758));
  AOI21_X1  g333(.A(KEYINPUT99), .B1(new_n758), .B2(new_n469), .ZN(new_n759));
  OAI221_X1 g334(.A(G2104), .B1(G116), .B2(new_n469), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G2067), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n751), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n541), .A2(G16), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n710), .A2(G21), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n765), .B1(G1966), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  NOR2_X1   g346(.A1(G171), .A2(new_n710), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G5), .B2(new_n710), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n752), .B1(new_n775), .B2(G34), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(KEYINPUT101), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(KEYINPUT101), .B2(new_n777), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G160), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT102), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n774), .B1(new_n771), .B2(new_n773), .C1(G2084), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n611), .B2(G16), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT97), .B(G1348), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n752), .A2(G33), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n482), .A2(G139), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT100), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n469), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n787), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n797), .A2(G2072), .B1(G2084), .B2(new_n781), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n752), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n752), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT29), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G2090), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n796), .A2(new_n442), .B1(new_n801), .B2(G2090), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n786), .A2(new_n798), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n710), .A2(G20), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT23), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(G164), .A2(G29), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G27), .B2(G29), .ZN(new_n811));
  AOI22_X1  g386(.A1(G1956), .A2(new_n809), .B1(new_n811), .B2(new_n443), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n443), .B2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n752), .A2(G32), .ZN(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT26), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G129), .B2(new_n484), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n752), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT27), .B(G1996), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT31), .B(G11), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT30), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n825), .A2(G28), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n752), .B1(new_n825), .B2(G28), .ZN(new_n827));
  OAI221_X1 g402(.A(new_n824), .B1(new_n826), .B2(new_n827), .C1(new_n634), .C2(new_n752), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n769), .B2(G1966), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n749), .A2(new_n750), .B1(new_n763), .B2(new_n762), .ZN(new_n830));
  INV_X1    g405(.A(G1956), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n808), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n823), .A2(new_n829), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  OR4_X1    g408(.A1(new_n782), .A2(new_n804), .A3(new_n813), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n747), .A2(new_n834), .ZN(G311));
  OR2_X1    g410(.A1(new_n747), .A2(new_n834), .ZN(G150));
  NAND2_X1  g411(.A1(new_n611), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI22_X1  g415(.A1(new_n513), .A2(new_n839), .B1(new_n840), .B2(new_n527), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n539), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n543), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n558), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n558), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n838), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(G860), .B1(new_n841), .B2(new_n843), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT103), .ZN(G145));
  XOR2_X1   g430(.A(new_n507), .B(new_n761), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n795), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(new_n819), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n819), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n484), .A2(G130), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n469), .A2(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(G142), .B2(new_n482), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n625), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n736), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n858), .A2(new_n867), .A3(new_n859), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n634), .B(KEYINPUT104), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G162), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G160), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n858), .A2(new_n867), .A3(KEYINPUT105), .A4(new_n859), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n878), .A2(new_n869), .A3(new_n879), .A4(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(G299), .A2(KEYINPUT106), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n568), .A2(new_n572), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n611), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n603), .A2(new_n610), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(KEYINPUT106), .A3(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(KEYINPUT41), .B2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(new_n847), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n620), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n890), .B(KEYINPUT107), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G288), .ZN(new_n899));
  XNOR2_X1  g474(.A(G303), .B(G305), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  OR3_X1    g478(.A1(new_n898), .A2(KEYINPUT110), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT110), .B1(new_n898), .B2(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n898), .A2(new_n903), .A3(KEYINPUT111), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G868), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n844), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n844), .ZN(G331));
  NAND2_X1  g488(.A1(new_n890), .A2(KEYINPUT41), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n914), .B(KEYINPUT114), .C1(new_n890), .C2(new_n891), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n615), .A2(G171), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(new_n541), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n894), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(KEYINPUT112), .ZN(new_n919));
  NOR2_X1   g494(.A1(G286), .A2(G301), .ZN(new_n920));
  INV_X1    g495(.A(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n847), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n922), .A3(KEYINPUT112), .ZN(new_n923));
  OR3_X1    g498(.A1(new_n890), .A2(KEYINPUT114), .A3(new_n891), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n915), .A2(new_n919), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT115), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n922), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n897), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n890), .B(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n930), .A2(KEYINPUT115), .A3(new_n922), .A4(new_n918), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n901), .B(KEYINPUT113), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n919), .A2(new_n923), .ZN(new_n935));
  INV_X1    g510(.A(new_n890), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(new_n893), .B2(new_n927), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n937), .B2(new_n901), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n934), .A2(new_n938), .A3(KEYINPUT43), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n893), .A2(new_n927), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n890), .B1(new_n919), .B2(new_n923), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT43), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n934), .A2(new_n938), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n938), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n949), .ZN(G397));
  INV_X1    g525(.A(KEYINPUT116), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n495), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n484), .A2(G126), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n503), .A2(new_n505), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n498), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G160), .A2(G40), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n507), .B2(new_n952), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n475), .A2(new_n963), .A3(new_n480), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(KEYINPUT116), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n761), .B(new_n763), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n819), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n737), .A2(new_n740), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n737), .A2(new_n740), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n819), .B(G1996), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n966), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n979), .A2(new_n966), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  INV_X1    g559(.A(new_n978), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n976), .A2(new_n985), .B1(G2067), .B2(new_n761), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n966), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n974), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n507), .A2(new_n990), .A3(new_n952), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n964), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2090), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n960), .B1(new_n957), .B2(new_n958), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n995));
  AOI21_X1  g570(.A(G1971), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(G8), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G303), .A2(G8), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(G8), .C1(new_n993), .C2(new_n996), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n964), .A2(new_n507), .A3(new_n952), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n583), .A2(new_n589), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n585), .A2(new_n591), .ZN(new_n1009));
  INV_X1    g584(.A(G1981), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT118), .A4(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G305), .B2(G1981), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n583), .B(new_n589), .C1(new_n584), .C2(new_n527), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1011), .A2(new_n1013), .B1(G1981), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1007), .B1(new_n1015), .B2(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1015), .A2(new_n1022), .A3(KEYINPUT49), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1016), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1006), .B(G8), .C1(new_n1025), .C2(G288), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n716), .B2(G1976), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(KEYINPUT52), .B2(new_n1026), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n959), .A2(new_n443), .A3(new_n995), .A4(new_n964), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT126), .B(KEYINPUT53), .Z(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n992), .A2(new_n771), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n962), .B2(new_n960), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n498), .A2(new_n955), .A3(new_n954), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n1040), .B2(new_n496), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT120), .B(new_n964), .C1(new_n1041), .C2(KEYINPUT45), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(new_n1042), .A3(new_n995), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G301), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1005), .A2(new_n1032), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1042), .A3(new_n995), .ZN(new_n1048));
  INV_X1    g623(.A(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n992), .A2(G2084), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(G168), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(KEYINPUT125), .B2(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(G8), .A3(new_n541), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT62), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1055), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n1058), .A4(new_n1056), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1047), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1017), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1024), .B2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1070), .A2(new_n1007), .B1(new_n1031), .B2(new_n1004), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1057), .A2(G8), .A3(new_n615), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1005), .A2(new_n1032), .A3(new_n1073), .A4(KEYINPUT63), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1003), .A2(new_n1024), .A3(new_n1004), .A4(new_n1030), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n1072), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1071), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1067), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n994), .A2(new_n995), .A3(new_n1044), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1035), .A2(new_n1036), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1045), .A2(new_n1035), .A3(G301), .A4(new_n1036), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(KEYINPUT54), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1064), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1081), .A2(G171), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1046), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n959), .A2(new_n995), .A3(new_n964), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n994), .A2(KEYINPUT121), .A3(new_n995), .A4(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n568), .A2(new_n572), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n831), .B2(new_n992), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1100), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n992), .A2(new_n831), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1006), .A2(G2067), .ZN(new_n1106));
  INV_X1    g681(.A(G1348), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n992), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n888), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1006), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n964), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n995), .A2(new_n967), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(KEYINPUT122), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n959), .A2(new_n967), .A3(new_n995), .A4(new_n964), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n1117), .B2(new_n1112), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n558), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1121), .B(new_n558), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1102), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(new_n1105), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n888), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n888), .B1(new_n1108), .B2(KEYINPUT60), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1127), .A2(new_n1128), .B1(KEYINPUT60), .B2(new_n1108), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1123), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1102), .A2(KEYINPUT61), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1105), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1124), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1094), .A2(new_n1095), .B1(new_n831), .B2(new_n992), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1134), .B(KEYINPUT123), .C1(new_n1103), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1110), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1090), .B1(new_n1138), .B2(KEYINPUT124), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(new_n1110), .C1(new_n1130), .C2(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1079), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n979), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n598), .B(G1986), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n980), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n988), .B1(new_n1142), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g721(.A1(new_n684), .A2(G319), .A3(new_n685), .ZN(new_n1148));
  NOR2_X1   g722(.A1(G229), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g723(.A1(new_n882), .A2(new_n663), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g724(.A1(new_n938), .A2(new_n942), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n1151), .A2(KEYINPUT43), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n934), .A2(new_n938), .A3(new_n946), .ZN(new_n1153));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(G308));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  NAND4_X1  g729(.A1(new_n1155), .A2(new_n663), .A3(new_n882), .A4(new_n1149), .ZN(G225));
endmodule


