//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1032,
    new_n1033, new_n1034;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  XNOR2_X1  g001(.A(G141gat), .B(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n203), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n203), .A2(KEYINPUT77), .ZN(new_n210));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n205), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT76), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G155gat), .B2(G162gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(new_n204), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222));
  OR2_X1    g021(.A1(G113gat), .A2(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G113gat), .A2(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n228), .A3(new_n224), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n229), .B(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n221), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n220), .ZN(new_n235));
  INV_X1    g034(.A(new_n209), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT78), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT78), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT2), .B1(new_n203), .B2(KEYINPUT77), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n219), .B1(new_n239), .B2(new_n214), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n240), .B2(new_n209), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n242), .B2(new_n233), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n202), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n237), .A2(new_n241), .A3(KEYINPUT3), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n233), .B1(new_n221), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n234), .A2(KEYINPUT4), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n221), .A2(new_n233), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n250), .A2(new_n254), .A3(new_n244), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n247), .B2(new_n249), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n251), .A2(new_n257), .A3(new_n253), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT83), .ZN(new_n264));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n256), .A2(new_n270), .A3(new_n262), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT40), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n244), .B1(new_n259), .B2(new_n260), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT39), .B1(new_n243), .B2(new_n245), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n258), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n260), .A3(new_n250), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n245), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT39), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n273), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(KEYINPUT39), .C1(new_n245), .C2(new_n243), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT39), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n282), .A2(KEYINPUT40), .A3(new_n268), .A4(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n272), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT70), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n295), .B2(KEYINPUT69), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n287), .B(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT69), .B1(new_n299), .B2(new_n289), .ZN(new_n300));
  INV_X1    g099(.A(new_n295), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G226gat), .ZN(new_n303));
  INV_X1    g102(.A(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT27), .B1(new_n306), .B2(KEYINPUT65), .ZN(new_n307));
  INV_X1    g106(.A(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT27), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G183gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n307), .B(new_n308), .C1(KEYINPUT65), .C2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT27), .B(G183gat), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n308), .A2(KEYINPUT28), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n317), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT67), .B1(new_n320), .B2(KEYINPUT26), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n322), .A3(new_n318), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n315), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n329), .A2(G169gat), .A3(G176gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n316), .A2(KEYINPUT23), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n332), .B(new_n325), .C1(KEYINPUT64), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n317), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(KEYINPUT64), .B(new_n335), .C1(new_n336), .C2(new_n317), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n325), .B(new_n335), .C1(new_n336), .C2(new_n317), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT25), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n334), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n334), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n328), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n305), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n337), .A2(new_n338), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT25), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n341), .B1(KEYINPUT25), .B2(new_n340), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n339), .A3(new_n342), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n327), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n305), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n302), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n302), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n345), .A2(new_n305), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(KEYINPUT29), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n305), .ZN(new_n360));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  NAND4_X1  g162(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT30), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n363), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n356), .A2(new_n360), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n356), .B2(new_n360), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n360), .A3(new_n363), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n371), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n286), .B1(new_n366), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n374), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n364), .B(KEYINPUT74), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n371), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n286), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT81), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n221), .A2(new_n248), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n346), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n302), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n304), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n297), .C1(new_n300), .C2(new_n301), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n242), .B1(new_n397), .B2(new_n248), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n389), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n248), .ZN(new_n400));
  INV_X1    g199(.A(new_n242), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n394), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n391), .B2(new_n302), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n346), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n299), .B2(new_n295), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n288), .A2(new_n301), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT3), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n392), .B1(new_n409), .B2(new_n221), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n399), .A2(new_n405), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n388), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n411), .A2(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n405), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n403), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n419), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n413), .A2(new_n417), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n411), .A2(new_n412), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n388), .A3(new_n424), .A4(new_n416), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n356), .A2(new_n360), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n356), .A2(new_n360), .A3(new_n368), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n367), .B1(new_n429), .B2(KEYINPUT37), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n268), .B1(new_n256), .B2(new_n262), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT6), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n435), .B2(KEYINPUT6), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n356), .A2(new_n360), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n363), .B1(new_n440), .B2(new_n428), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n354), .B1(new_n353), .B2(new_n406), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n358), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n428), .B1(new_n443), .B2(new_n357), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n302), .B(new_n358), .C1(new_n359), .C2(new_n305), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n427), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n441), .A2(new_n446), .B1(new_n440), .B2(new_n363), .ZN(new_n447));
  INV_X1    g246(.A(new_n278), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n448), .A2(new_n261), .B1(new_n246), .B2(new_n255), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT6), .B1(new_n449), .B2(new_n268), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n272), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n434), .A2(new_n439), .A3(new_n447), .A4(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n379), .A2(new_n387), .A3(new_n426), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n377), .A2(new_n366), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n263), .A2(new_n269), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n426), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n345), .A2(new_n233), .ZN(new_n460));
  INV_X1    g259(.A(new_n233), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n353), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G227gat), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n304), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT34), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n469), .A3(new_n466), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G15gat), .B(G43gat), .Z(new_n474));
  XNOR2_X1  g273(.A(G71gat), .B(G99gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n468), .B(new_n470), .C1(new_n473), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n471), .B2(new_n472), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n469), .B1(new_n463), .B2(new_n466), .ZN(new_n480));
  AOI211_X1 g279(.A(KEYINPUT34), .B(new_n465), .C1(new_n460), .C2(new_n462), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n471), .A2(KEYINPUT32), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n484), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n478), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(KEYINPUT36), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n478), .A2(new_n482), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n478), .B2(new_n482), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n458), .A2(new_n459), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n454), .A2(new_n494), .A3(new_n426), .A4(new_n457), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT35), .B1(new_n439), .B2(new_n451), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(new_n454), .A3(new_n494), .A4(new_n426), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n453), .A2(new_n493), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n502), .B(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT12), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT16), .ZN(new_n511));
  NAND2_X1  g310(.A1(G15gat), .A2(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(G15gat), .A2(G22gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G15gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n412), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(new_n510), .A3(new_n512), .ZN(new_n518));
  AOI211_X1 g317(.A(KEYINPUT87), .B(G8gat), .C1(new_n515), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n515), .A2(new_n518), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(G43gat), .A2(G50gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NAND2_X1  g328(.A1(G43gat), .A2(G50gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G29gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(G29gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n530), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT15), .B1(new_n540), .B2(new_n527), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n531), .A2(new_n541), .A3(new_n537), .A4(new_n538), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n526), .A2(KEYINPUT88), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT88), .B1(new_n526), .B2(new_n545), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n546), .A2(new_n547), .B1(new_n545), .B2(new_n526), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT13), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n552));
  INV_X1    g351(.A(new_n545), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n515), .A2(new_n518), .A3(new_n523), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n520), .A3(new_n521), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n524), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n526), .A2(new_n545), .A3(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n543), .A2(KEYINPUT17), .A3(new_n544), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n559), .A2(KEYINPUT18), .A3(new_n549), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n551), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n563), .B(new_n549), .C1(new_n546), .C2(new_n547), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n565), .B1(new_n551), .B2(new_n564), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n509), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n506), .A2(new_n508), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n569), .A2(new_n551), .A3(new_n564), .A4(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT90), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n509), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n577), .A2(KEYINPUT90), .A3(new_n551), .A4(new_n564), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n499), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G71gat), .ZN(new_n586));
  INV_X1    g385(.A(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n585), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n589), .B(new_n588), .C1(new_n584), .C2(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n556), .B1(new_n583), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT92), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT91), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n597), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n595), .A2(new_n583), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n602), .B(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT8), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(G99gat), .B2(G106gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT93), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT8), .ZN(new_n617));
  OR2_X1    g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n611), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n610), .B(new_n626), .C1(new_n615), .C2(new_n620), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n609), .B1(new_n631), .B2(new_n553), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n561), .A2(new_n562), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n630), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT94), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n632), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n632), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641));
  INV_X1    g440(.A(G232gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n642), .B2(new_n304), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n640), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n637), .B2(new_n638), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n608), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n595), .B1(new_n628), .B2(new_n629), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n617), .A2(new_n619), .A3(new_n618), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n619), .B1(new_n617), .B2(new_n618), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n627), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n610), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n593), .A2(new_n594), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n621), .A2(new_n611), .A3(new_n627), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n650), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n650), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n651), .A2(new_n663), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n656), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G120gat), .B(G148gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(G176gat), .B(G204gat), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n667), .B(new_n668), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n661), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n666), .B2(new_n659), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n649), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n582), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT96), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n582), .A2(KEYINPUT96), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT6), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT80), .B1(new_n455), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT6), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n456), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g485(.A(new_n454), .B1(new_n678), .B2(new_n679), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n521), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n689), .B2(new_n691), .ZN(G1325gat));
  NAND3_X1  g492(.A1(new_n680), .A2(new_n516), .A3(new_n494), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n492), .A2(new_n488), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n678), .B2(new_n679), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(new_n516), .ZN(G1326gat));
  INV_X1    g496(.A(KEYINPUT97), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n680), .B2(new_n459), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT97), .B(new_n426), .C1(new_n678), .C2(new_n679), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n699), .B2(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n582), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n608), .A2(new_n674), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n648), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n535), .A3(new_n684), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n499), .B2(new_n648), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n648), .A2(KEYINPUT101), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n646), .B2(new_n647), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT100), .B(KEYINPUT44), .Z(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n715), .B1(new_n499), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n684), .A2(new_n385), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n695), .B1(new_n725), .B2(new_n426), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n452), .A2(new_n426), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n386), .B1(new_n385), .B2(new_n286), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(new_n387), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n496), .A2(new_n498), .ZN(new_n731));
  OAI211_X1 g530(.A(KEYINPUT102), .B(new_n722), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n714), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT98), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n572), .A2(new_n579), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n572), .B2(new_n579), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n707), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT99), .Z(new_n739));
  NAND3_X1  g538(.A1(new_n733), .A2(new_n684), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n535), .B1(new_n740), .B2(KEYINPUT103), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(KEYINPUT103), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n713), .A2(new_n742), .ZN(G1328gat));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n711), .A2(new_n532), .A3(new_n385), .A4(new_n745), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n744), .A2(KEYINPUT104), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n733), .A2(new_n385), .A3(new_n739), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n532), .B2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(new_n695), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n751), .A3(new_n739), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n751), .A4(new_n739), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(G43gat), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n494), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n582), .A2(new_n709), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n752), .A2(G43gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n759), .B1(new_n752), .B2(G43gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(KEYINPUT105), .A3(KEYINPUT47), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(G1330gat));
  NAND4_X1  g568(.A1(new_n733), .A2(G50gat), .A3(new_n459), .A4(new_n739), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n706), .A2(new_n426), .A3(new_n710), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(G50gat), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g572(.A1(new_n737), .A2(new_n649), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n674), .ZN(new_n775));
  XOR2_X1   g574(.A(new_n775), .B(KEYINPUT107), .Z(new_n776));
  INV_X1    g575(.A(new_n499), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n684), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g580(.A(new_n454), .B(new_n778), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  NOR3_X1   g583(.A1(new_n778), .A2(G71gat), .A3(new_n757), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n751), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(G71gat), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g587(.A1(new_n778), .A2(new_n426), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n587), .ZN(G1335gat));
  NOR4_X1   g589(.A1(new_n499), .A2(new_n608), .A3(new_n648), .A4(new_n737), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(KEYINPUT51), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(KEYINPUT51), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n457), .A2(G85gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n674), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n737), .A2(new_n608), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n674), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n733), .A2(new_n684), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G85gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1336gat));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n454), .A2(G92gat), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n674), .B(new_n804), .C1(new_n792), .C2(new_n793), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n733), .A2(new_n385), .A3(new_n799), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n803), .B(new_n805), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(G92gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(G1337gat));
  NOR2_X1   g614(.A1(new_n757), .A2(G99gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n674), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n733), .A2(new_n751), .A3(new_n799), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G99gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1338gat));
  INV_X1    g619(.A(new_n674), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n426), .A2(G106gat), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT109), .Z(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n792), .B2(new_n793), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n733), .A2(new_n459), .A3(new_n799), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g627(.A(new_n608), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n664), .A2(new_n665), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n650), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n664), .A2(new_n662), .A3(new_n665), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT110), .B(new_n669), .C1(new_n666), .C2(new_n832), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n833), .A2(new_n832), .A3(new_n650), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n670), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT111), .B(new_n836), .C1(new_n837), .C2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  AOI211_X1 g641(.A(KEYINPUT54), .B(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT110), .B1(new_n843), .B2(new_n669), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n838), .A3(new_n670), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT111), .B1(new_n846), .B2(new_n836), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n844), .A2(new_n845), .B1(new_n835), .B2(new_n834), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n672), .B1(new_n849), .B2(KEYINPUT55), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n830), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n836), .B1(new_n837), .B2(new_n840), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n841), .ZN(new_n855));
  INV_X1    g654(.A(new_n672), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n835), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(new_n831), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT112), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n851), .A2(new_n737), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n548), .A2(new_n550), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n549), .B1(new_n559), .B2(new_n563), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n504), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT113), .Z(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n674), .A3(new_n579), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n719), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n579), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n719), .A3(new_n860), .A4(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n829), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n774), .A2(new_n821), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n457), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n494), .A2(new_n426), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n385), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(G113gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n581), .ZN(new_n878));
  INV_X1    g677(.A(new_n876), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n737), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n877), .B2(new_n880), .ZN(G1340gat));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n674), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g682(.A1(new_n876), .A2(new_n829), .ZN(new_n884));
  XNOR2_X1  g683(.A(KEYINPUT114), .B(G127gat), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n884), .B(new_n885), .ZN(G1342gat));
  NOR2_X1   g685(.A1(new_n385), .A2(new_n648), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT115), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(G134gat), .A3(new_n874), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT56), .Z(new_n891));
  OAI21_X1  g690(.A(G134gat), .B1(new_n876), .B2(new_n648), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n872), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n459), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n695), .A2(new_n684), .A3(new_n454), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n855), .A2(new_n859), .A3(new_n580), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n866), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n648), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n608), .B1(new_n869), .B2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n872), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n459), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n897), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n580), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n896), .A2(new_n907), .A3(new_n904), .A4(new_n580), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(G141gat), .A3(new_n908), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n426), .B(new_n897), .C1(new_n871), .C2(new_n872), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n581), .A2(G141gat), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT58), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n904), .ZN(new_n917));
  INV_X1    g716(.A(new_n737), .ZN(new_n918));
  OAI21_X1  g717(.A(G141gat), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n910), .A2(new_n911), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT58), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n914), .A2(new_n916), .A3(new_n922), .ZN(G1344gat));
  INV_X1    g722(.A(G148gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n910), .A2(new_n924), .A3(new_n674), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n675), .A2(new_n581), .ZN(new_n927));
  INV_X1    g726(.A(new_n648), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n868), .A2(new_n928), .A3(new_n855), .A4(new_n859), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n900), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n930), .B2(new_n608), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT57), .B1(new_n931), .B2(new_n459), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n861), .A2(new_n866), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n720), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n608), .B1(new_n934), .B2(new_n869), .ZN(new_n935));
  OAI211_X1 g734(.A(KEYINPUT57), .B(new_n459), .C1(new_n935), .C2(new_n902), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n932), .B1(new_n936), .B2(KEYINPUT119), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n895), .B(new_n426), .C1(new_n871), .C2(new_n872), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n821), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n897), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n926), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n924), .A2(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n917), .B2(new_n821), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n925), .B1(new_n944), .B2(new_n948), .ZN(G1345gat));
  OAI21_X1  g748(.A(G155gat), .B1(new_n917), .B2(new_n829), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n910), .A2(new_n206), .A3(new_n608), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT120), .Z(G1346gat));
  NOR4_X1   g752(.A1(new_n888), .A2(G162gat), .A3(new_n457), .A4(new_n751), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n894), .A2(new_n954), .A3(new_n459), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT121), .Z(new_n956));
  OAI21_X1  g755(.A(G162gat), .B1(new_n917), .B2(new_n720), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1347gat));
  AOI21_X1  g757(.A(new_n684), .B1(new_n871), .B2(new_n872), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n874), .A2(new_n454), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(G169gat), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n961), .A2(new_n962), .A3(new_n581), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n894), .A2(new_n457), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n960), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT123), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n971), .A3(new_n960), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n737), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n963), .B1(new_n973), .B2(new_n962), .ZN(G1348gat));
  NOR2_X1   g773(.A1(new_n821), .A2(G176gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G176gat), .B1(new_n961), .B2(new_n821), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1349gat));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n608), .A2(new_n313), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n968), .A2(new_n960), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G183gat), .B1(new_n961), .B2(new_n829), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  NOR2_X1   g786(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n987), .ZN(new_n989));
  AOI211_X1 g788(.A(new_n980), .B(new_n989), .C1(new_n983), .C2(new_n984), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n988), .A2(new_n990), .ZN(G1350gat));
  NAND4_X1  g790(.A1(new_n970), .A2(new_n308), .A3(new_n719), .A4(new_n972), .ZN(new_n992));
  OAI21_X1  g791(.A(G190gat), .B1(new_n961), .B2(new_n648), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1351gat));
  NOR3_X1   g794(.A1(new_n751), .A2(new_n454), .A3(new_n426), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n968), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(G197gat), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n737), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n751), .A2(new_n684), .A3(new_n454), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n931), .A2(new_n459), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(new_n895), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1002), .B1(new_n938), .B2(new_n939), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n580), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G197gat), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n999), .B1(new_n1008), .B2(new_n1009), .ZN(G1352gat));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g810(.A(G204gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1012), .B1(new_n941), .B2(new_n1000), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT62), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n821), .A2(G204gat), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n968), .A2(new_n1014), .A3(new_n996), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT122), .B1(new_n894), .B2(new_n457), .ZN(new_n1017));
  AOI211_X1 g816(.A(new_n965), .B(new_n684), .C1(new_n871), .C2(new_n872), .ZN(new_n1018));
  OAI211_X1 g817(.A(new_n996), .B(new_n1015), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1011), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g821(.A(new_n674), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1023), .A2(G204gat), .ZN(new_n1024));
  NAND4_X1  g823(.A1(new_n1024), .A2(KEYINPUT127), .A3(new_n1020), .A4(new_n1016), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1022), .A2(new_n1025), .ZN(G1353gat));
  NAND3_X1  g825(.A1(new_n997), .A2(new_n292), .A3(new_n608), .ZN(new_n1027));
  OAI211_X1 g826(.A(new_n608), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n1028), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1029));
  AOI21_X1  g828(.A(KEYINPUT63), .B1(new_n1028), .B2(G211gat), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G1354gat));
  NAND3_X1  g830(.A1(new_n997), .A2(new_n293), .A3(new_n719), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n937), .A2(new_n940), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1033), .A2(new_n928), .A3(new_n1000), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1032), .B1(new_n1034), .B2(new_n293), .ZN(G1355gat));
endmodule


