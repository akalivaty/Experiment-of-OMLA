//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT3), .A3(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n189), .B1(new_n197), .B2(G101), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  AND4_X1   g014(.A1(new_n199), .A2(new_n195), .A3(new_n200), .A4(new_n196), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n192), .A2(new_n194), .B1(new_n191), .B2(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n199), .B1(new_n202), .B2(new_n200), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n198), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT70), .A2(G116), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT70), .A2(G116), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G119), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT2), .B(G113), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n211), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n207), .A3(new_n209), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n200), .B1(new_n195), .B2(new_n196), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n212), .A2(new_n214), .B1(new_n215), .B2(new_n189), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n204), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n195), .A2(new_n200), .A3(new_n196), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT76), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n202), .A2(new_n199), .A3(new_n200), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n196), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n191), .A2(KEYINPUT77), .A3(G107), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n223), .B(new_n224), .C1(new_n191), .C2(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n207), .A2(KEYINPUT5), .A3(new_n209), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n227), .B(G113), .C1(KEYINPUT5), .C2(new_n209), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n221), .A2(new_n214), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G110), .B(G122), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT81), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n217), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT6), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n217), .B2(new_n229), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G224), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G953), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  INV_X1    g052(.A(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(G128), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT64), .B1(new_n239), .B2(G143), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G128), .A4(new_n240), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n245), .A2(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n243), .B2(new_n246), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT69), .A3(new_n248), .A4(G128), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n242), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G125), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT0), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n238), .B2(new_n258), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n258), .B(new_n252), .C1(new_n243), .C2(new_n246), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT0), .B1(new_n238), .B2(G128), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n237), .B1(new_n256), .B2(new_n264), .ZN(new_n265));
  OAI221_X1 g079(.A(new_n263), .B1(new_n236), .B2(G953), .C1(new_n255), .C2(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT6), .B(new_n231), .C1(new_n217), .C2(new_n229), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n235), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n231), .B(KEYINPUT8), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n226), .B1(new_n201), .B2(new_n203), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n228), .A2(new_n214), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n221), .A2(new_n226), .B1(new_n228), .B2(new_n214), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT7), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n237), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n256), .B2(new_n264), .ZN(new_n278));
  OAI221_X1 g092(.A(new_n263), .B1(new_n276), .B2(new_n237), .C1(new_n255), .C2(G125), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(new_n278), .A3(new_n232), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n188), .B1(new_n269), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n282), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n217), .A2(new_n229), .ZN(new_n285));
  INV_X1    g099(.A(new_n231), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT6), .A3(new_n232), .ZN(new_n288));
  INV_X1    g102(.A(new_n268), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n265), .A4(new_n266), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n284), .A2(new_n290), .A3(new_n187), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT82), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT82), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  XNOR2_X1  g111(.A(G128), .B(G143), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n205), .A2(G122), .A3(new_n206), .ZN(new_n301));
  INV_X1    g115(.A(G122), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G116), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT14), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT14), .ZN(new_n306));
  OAI21_X1  g120(.A(G107), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  OAI221_X1 g121(.A(new_n300), .B1(G107), .B2(new_n304), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT13), .B1(new_n258), .B2(G143), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n299), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n298), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n193), .B1(new_n301), .B2(new_n303), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n304), .A2(G107), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  INV_X1    g130(.A(G217), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n316), .A2(new_n317), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n308), .A2(new_n314), .A3(new_n318), .ZN(new_n321));
  AOI21_X1  g135(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G478), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT15), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n325), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT87), .B(G952), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G953), .ZN(new_n330));
  NAND2_X1  g144(.A1(G234), .A2(G237), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT88), .Z(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(G902), .A3(G953), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT21), .B(G898), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G475), .ZN(new_n339));
  NOR2_X1   g153(.A1(G237), .A2(G953), .ZN(new_n340));
  AOI21_X1  g154(.A(G143), .B1(new_n340), .B2(G214), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(G143), .A3(G214), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT18), .A2(G131), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  OAI211_X1 g160(.A(KEYINPUT18), .B(G131), .C1(new_n346), .C2(new_n341), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(new_n239), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n239), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(KEYINPUT83), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n348), .A2(new_n352), .A3(new_n239), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n345), .B(new_n347), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n356), .A2(KEYINPUT16), .ZN(new_n357));
  INV_X1    g171(.A(G125), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G140), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(KEYINPUT16), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(G146), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(G146), .B1(new_n357), .B2(new_n360), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT17), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT66), .B(G131), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n346), .B2(new_n341), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n364), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n342), .A2(new_n366), .A3(new_n343), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(KEYINPUT17), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n354), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(G113), .B(G122), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n191), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n375), .B(new_n354), .C1(new_n369), .C2(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n339), .B1(new_n379), .B2(new_n281), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n348), .A2(KEYINPUT84), .A3(KEYINPUT19), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT19), .B1(new_n348), .B2(KEYINPUT84), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n239), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n371), .A3(new_n361), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n354), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n376), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT85), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n388), .A3(new_n376), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n378), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G475), .A2(G902), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT86), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n380), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n378), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n388), .B1(new_n385), .B2(new_n376), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n390), .A2(KEYINPUT86), .A3(new_n391), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT20), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n338), .A2(new_n394), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n338), .A2(new_n394), .A3(KEYINPUT89), .A4(new_n401), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n295), .A2(new_n297), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n299), .B2(G137), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT67), .ZN(new_n411));
  INV_X1    g225(.A(G137), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(G134), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n299), .A2(KEYINPUT67), .A3(G137), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(G134), .ZN(new_n416));
  OR2_X1    g230(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n417), .B2(new_n409), .ZN(new_n418));
  OAI21_X1  g232(.A(G131), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT68), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n412), .A2(G134), .ZN(new_n422));
  AOI22_X1  g236(.A1(KEYINPUT67), .A2(new_n422), .B1(new_n416), .B2(new_n409), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n299), .A2(G137), .ZN(new_n424));
  INV_X1    g238(.A(new_n409), .ZN(new_n425));
  NOR2_X1   g239(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n423), .A2(new_n427), .A3(new_n366), .A4(new_n413), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT68), .B(G131), .C1(new_n415), .C2(new_n418), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n421), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT10), .B(new_n226), .C1(new_n201), .C2(new_n203), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n215), .A2(new_n189), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n262), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT4), .B1(new_n202), .B2(new_n200), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n219), .B2(new_n220), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n255), .A2(new_n432), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n251), .A2(new_n254), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n248), .B1(G143), .B2(new_n239), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n258), .B1(new_n441), .B2(KEYINPUT78), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n241), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n253), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n219), .A2(new_n220), .B1(G101), .B2(new_n225), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT10), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n445), .B1(new_n251), .B2(new_n254), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n439), .B(new_n450), .C1(new_n452), .C2(new_n271), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n431), .B(new_n438), .C1(new_n451), .C2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n456));
  INV_X1    g270(.A(new_n242), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n440), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n448), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n452), .A2(new_n271), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT12), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n456), .B(new_n463), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  INV_X1    g280(.A(G953), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G227), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n466), .B(new_n468), .Z(new_n469));
  OAI21_X1  g283(.A(new_n450), .B1(new_n452), .B2(new_n271), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT79), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n437), .B1(new_n471), .B2(new_n453), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n469), .B1(new_n472), .B2(new_n431), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n438), .B1(new_n451), .B2(new_n454), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n430), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n465), .A2(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G469), .B1(new_n476), .B2(G902), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n472), .A2(new_n431), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n430), .B(new_n437), .C1(new_n471), .C2(new_n453), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n469), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n455), .A2(new_n481), .A3(new_n462), .A4(new_n464), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G469), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n281), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n408), .B1(new_n477), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n406), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n208), .B2(G128), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n490), .B(new_n491), .C1(G119), .C2(new_n258), .ZN(new_n492));
  XNOR2_X1  g306(.A(G119), .B(G128), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT24), .B(G110), .Z(new_n494));
  OAI22_X1  g308(.A1(new_n492), .A2(G110), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n361), .A3(new_n350), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(G110), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n494), .A2(KEYINPUT74), .A3(new_n493), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT74), .B1(new_n494), .B2(new_n493), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n496), .B1(new_n364), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n467), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n496), .B(new_n504), .C1(new_n364), .C2(new_n500), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n281), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n506), .A2(KEYINPUT25), .A3(new_n281), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n317), .B1(G234), .B2(new_n281), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n488), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n513), .ZN(new_n515));
  AOI211_X1 g329(.A(KEYINPUT75), .B(new_n515), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n506), .A2(new_n507), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n513), .A2(G902), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G472), .ZN(new_n523));
  INV_X1    g337(.A(new_n259), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n253), .A2(G128), .ZN(new_n525));
  INV_X1    g339(.A(new_n261), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n429), .A2(new_n428), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n421), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n422), .B2(new_n424), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n428), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n440), .B2(new_n457), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n212), .A2(new_n214), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT30), .B1(new_n529), .B2(new_n532), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n419), .A2(new_n420), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n429), .A2(new_n428), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n262), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n538), .B(new_n539), .C1(new_n255), .C2(new_n531), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n534), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n340), .A2(G210), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n543), .B(KEYINPUT27), .Z(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n546), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT28), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n533), .B1(new_n529), .B2(new_n532), .ZN(new_n550));
  INV_X1    g364(.A(new_n533), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n538), .B(new_n551), .C1(new_n255), .C2(new_n531), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n549), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n529), .A2(new_n532), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT28), .B1(new_n554), .B2(new_n551), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n548), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n547), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT72), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  INV_X1    g372(.A(new_n531), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n458), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n551), .B1(new_n560), .B2(new_n538), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT28), .B1(new_n534), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n548), .A2(KEYINPUT29), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n281), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n567), .B2(KEYINPUT73), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n569), .A3(new_n281), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n523), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n542), .B2(new_n548), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n551), .B1(new_n535), .B2(new_n540), .ZN(new_n576));
  NOR4_X1   g390(.A1(new_n576), .A2(KEYINPUT31), .A3(new_n534), .A4(new_n546), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n552), .A2(new_n549), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n548), .B1(new_n562), .B2(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(G472), .A2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n573), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n542), .A2(new_n548), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT31), .ZN(new_n585));
  INV_X1    g399(.A(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n542), .A2(new_n574), .A3(new_n548), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT32), .A3(new_n581), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n522), .B1(new_n571), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n487), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT90), .B(G101), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G3));
  AND2_X1   g408(.A1(new_n486), .A2(new_n522), .ZN(new_n595));
  INV_X1    g409(.A(new_n293), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n187), .B1(new_n284), .B2(new_n290), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n597), .B2(KEYINPUT91), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n283), .A2(new_n291), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n394), .A2(new_n401), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT93), .B(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n322), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n320), .A2(new_n321), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n606), .A2(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n320), .A2(KEYINPUT92), .A3(new_n606), .A4(new_n321), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n323), .A2(G902), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n604), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n602), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n601), .A2(new_n615), .A3(new_n337), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n523), .B1(new_n588), .B2(new_n281), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n588), .B2(new_n581), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n595), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT94), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT34), .B(G104), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n337), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n394), .A2(new_n401), .A3(new_n623), .A4(new_n328), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n601), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n595), .A2(new_n618), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n501), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n519), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n517), .A2(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(G469), .B(G902), .C1(new_n480), .C2(new_n482), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n462), .A2(new_n464), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n469), .B1(new_n634), .B2(new_n479), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n473), .A2(new_n475), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(G469), .ZN(new_n637));
  NAND2_X1  g451(.A1(G469), .A2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n407), .B(new_n632), .C1(new_n633), .C2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n406), .A2(new_n641), .A3(new_n618), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  NOR2_X1   g458(.A1(new_n571), .A2(new_n590), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n598), .A2(new_n600), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n486), .A2(new_n646), .A3(new_n632), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n334), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n333), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n394), .A2(new_n401), .A3(new_n328), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n645), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n258), .ZN(G30));
  XNOR2_X1  g472(.A(new_n292), .B(KEYINPUT38), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n328), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n394), .B2(new_n401), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR4_X1   g477(.A1(new_n660), .A2(new_n596), .A3(new_n632), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n650), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n486), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n542), .A2(new_n546), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n550), .A2(new_n552), .A3(new_n546), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n281), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n583), .A2(new_n589), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n664), .A2(new_n667), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  AND3_X1   g489(.A1(new_n566), .A2(new_n569), .A3(new_n281), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n569), .B1(new_n566), .B2(new_n281), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n677), .A3(new_n557), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n589), .B(new_n583), .C1(new_n678), .C2(new_n523), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n640), .A2(new_n601), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n613), .B1(new_n394), .B2(new_n401), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n651), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AOI21_X1  g499(.A(new_n481), .B1(new_n475), .B2(new_n455), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n455), .A2(new_n481), .A3(new_n462), .A4(new_n464), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n281), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n407), .A3(new_n485), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT96), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n689), .A2(KEYINPUT96), .A3(new_n407), .A4(new_n485), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n616), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n591), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT41), .B(G113), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n625), .A3(new_n693), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n591), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(G116), .Z(G18));
  NOR2_X1   g514(.A1(new_n690), .A2(new_n601), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n630), .A2(new_n519), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n514), .A2(new_n516), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(new_n404), .B2(new_n405), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n645), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n208), .ZN(G21));
  AND4_X1   g521(.A1(new_n623), .A2(new_n662), .A3(new_n598), .A4(new_n600), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n692), .A2(new_n693), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT97), .B(G472), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n580), .B2(G902), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n558), .A2(new_n564), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n585), .B(new_n587), .C1(new_n712), .C2(new_n548), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n711), .A2(KEYINPUT98), .B1(new_n581), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n710), .C1(new_n580), .C2(G902), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n522), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n302), .ZN(G24));
  NAND2_X1  g533(.A1(new_n701), .A2(new_n683), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n713), .A2(new_n581), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n632), .A3(new_n716), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n714), .A2(KEYINPUT99), .A3(new_n632), .A4(new_n716), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n358), .ZN(G27));
  NAND2_X1  g542(.A1(new_n568), .A2(new_n570), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G472), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT32), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n580), .B2(new_n582), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n589), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n734), .B(new_n407), .C1(new_n633), .C2(new_n639), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n682), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n522), .A4(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n679), .A2(new_n736), .A3(KEYINPUT100), .A4(new_n522), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n583), .A2(new_n589), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n521), .B1(new_n730), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT100), .B1(new_n742), .B2(new_n736), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n737), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND4_X1  g559(.A1(new_n654), .A2(new_n486), .A3(new_n655), .A4(new_n734), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n591), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n299), .ZN(G36));
  AND2_X1   g562(.A1(new_n394), .A2(new_n401), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n614), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n632), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n618), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT103), .Z(new_n756));
  NAND2_X1  g570(.A1(new_n635), .A2(new_n636), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n484), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n638), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT101), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n633), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n407), .ZN(new_n766));
  INV_X1    g580(.A(new_n665), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n766), .A2(KEYINPUT102), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT102), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  INV_X1    g583(.A(new_n734), .ZN(new_n770));
  OR3_X1    g584(.A1(new_n754), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT104), .B1(new_n754), .B2(KEYINPUT44), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n756), .A2(new_n768), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  XNOR2_X1  g589(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n766), .B(new_n777), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n679), .A2(new_n522), .A3(new_n682), .A4(new_n770), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(KEYINPUT106), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(new_n333), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n752), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n690), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n734), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n733), .A2(new_n522), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n793), .B(KEYINPUT48), .Z(new_n794));
  OR2_X1    g608(.A1(new_n787), .A2(new_n717), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n601), .A3(new_n690), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n789), .A2(new_n521), .A3(new_n333), .A4(new_n673), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n681), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n330), .B(KEYINPUT119), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n794), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n689), .A2(new_n485), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n408), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n778), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n795), .A2(new_n770), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n660), .A2(new_n596), .A3(new_n788), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n795), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(new_n810), .B2(KEYINPUT116), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n725), .A2(new_n726), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n790), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT117), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n602), .A2(new_n614), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n797), .B2(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT50), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n800), .B1(new_n808), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT118), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n816), .A2(new_n826), .A3(new_n821), .A4(new_n822), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n825), .B(new_n827), .C1(new_n805), .C2(new_n807), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n717), .A2(new_n709), .B1(new_n698), .B2(new_n591), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n591), .B1(new_n694), .B2(new_n487), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n295), .A2(new_n297), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n749), .A2(new_n328), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n337), .B1(new_n835), .B2(new_n615), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n595), .A2(new_n834), .A3(new_n618), .A4(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n837), .B(new_n642), .C1(new_n645), .C2(new_n705), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n661), .A2(new_n651), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n703), .A2(new_n602), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n486), .A2(new_n841), .A3(new_n734), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n591), .A2(new_n746), .B1(new_n645), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n817), .B2(new_n736), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n744), .A2(new_n833), .A3(new_n839), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT109), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n838), .A2(new_n831), .A3(new_n832), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n744), .A4(new_n844), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n720), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n657), .B1(new_n817), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n632), .B2(new_n650), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n703), .A2(KEYINPUT111), .A3(new_n651), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n601), .A2(new_n663), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n673), .A4(new_n486), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n684), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT112), .B1(new_n852), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n727), .A2(new_n859), .A3(new_n862), .A4(new_n657), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n861), .B2(new_n863), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n850), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n845), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n852), .A2(new_n860), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT52), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT53), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n846), .A2(KEYINPUT110), .A3(new_n849), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT110), .B1(new_n846), .B2(new_n849), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n867), .A2(new_n873), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n880), .A2(KEYINPUT53), .B1(new_n869), .B2(new_n868), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n876), .B1(new_n881), .B2(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n830), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n750), .A2(new_n521), .A3(new_n596), .A4(new_n408), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n801), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT107), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n659), .B1(new_n886), .B2(new_n801), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n741), .A3(new_n672), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT108), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n884), .A2(new_n891), .ZN(G75));
  INV_X1    g706(.A(new_n874), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n869), .B2(new_n868), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n281), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n235), .A2(new_n268), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n267), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n467), .A2(G952), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G51));
  XOR2_X1   g718(.A(new_n638), .B(KEYINPUT57), .Z(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n894), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n876), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT120), .B(new_n905), .C1(new_n876), .C2(new_n907), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n483), .A3(new_n911), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n894), .A2(new_n281), .A3(new_n760), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n903), .B1(new_n912), .B2(new_n913), .ZN(G54));
  NAND3_X1  g728(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n390), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n903), .ZN(G60));
  INV_X1    g733(.A(new_n611), .ZN(new_n920));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  OR2_X1    g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n894), .A2(new_n906), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n903), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n920), .B1(new_n882), .B2(new_n922), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n926), .B2(new_n903), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n869), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n846), .A2(new_n849), .B1(new_n864), .B2(KEYINPUT52), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n867), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n630), .B(new_n933), .C1(new_n936), .C2(new_n893), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  INV_X1    g752(.A(new_n903), .ZN(new_n939));
  INV_X1    g753(.A(new_n518), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n894), .B2(new_n932), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n938), .A2(KEYINPUT124), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n939), .A4(new_n937), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n937), .A2(KEYINPUT122), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n875), .A2(new_n948), .A3(new_n630), .A4(new_n933), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n947), .A2(new_n939), .A3(new_n949), .A4(new_n941), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT123), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(G66));
  OAI21_X1  g768(.A(G953), .B1(new_n335), .B2(new_n236), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n847), .B2(G953), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n235), .A2(new_n268), .B1(G898), .B2(new_n467), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  AOI21_X1  g772(.A(new_n681), .B1(new_n749), .B2(new_n328), .ZN(new_n959));
  OR4_X1    g773(.A1(new_n591), .A2(new_n666), .A3(new_n959), .A4(new_n770), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n852), .A2(new_n684), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n674), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NAND4_X1  g777(.A1(new_n784), .A2(new_n774), .A3(new_n960), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n467), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n381), .A2(new_n382), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n541), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(G900), .B2(G953), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n768), .A2(new_n857), .A3(new_n792), .A4(new_n769), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n774), .A2(new_n961), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n744), .B1(new_n591), .B2(new_n746), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT126), .Z(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(new_n784), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n974), .B2(G953), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n467), .B1(G227), .B2(G900), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n976), .B(new_n979), .ZN(G72));
  NAND2_X1  g794(.A1(G472), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT63), .Z(new_n982));
  INV_X1    g796(.A(new_n847), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n964), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n669), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n974), .B2(new_n983), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n547), .B(KEYINPUT127), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n669), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n881), .A2(new_n547), .A3(new_n989), .A4(new_n982), .ZN(new_n990));
  AND4_X1   g804(.A1(new_n939), .A2(new_n985), .A3(new_n988), .A4(new_n990), .ZN(G57));
endmodule


