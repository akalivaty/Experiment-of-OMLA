//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n203), .B2(new_n202), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT93), .B(G8gat), .Z(new_n206));
  AOI21_X1  g005(.A(KEYINPUT94), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(KEYINPUT94), .A3(new_n206), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(new_n205), .ZN(new_n210));
  AOI21_X1  g009(.A(G64gat), .B1(KEYINPUT98), .B2(G57gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT97), .A2(KEYINPUT98), .A3(G57gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT97), .B2(G57gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n213), .B2(G64gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT99), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT9), .ZN(new_n216));
  INV_X1    g015(.A(G71gat), .ZN(new_n217));
  INV_X1    g016(.A(G78gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G71gat), .B(G78gat), .Z(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n215), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n221), .A2(KEYINPUT96), .ZN(new_n223));
  OR2_X1    g022(.A1(G57gat), .A2(G64gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(G57gat), .A2(G64gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n221), .A2(KEYINPUT96), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  AOI211_X1 g028(.A(new_n207), .B(new_n210), .C1(new_n229), .C2(KEYINPUT21), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G155gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n229), .A2(KEYINPUT21), .ZN(new_n235));
  NAND2_X1  g034(.A1(G231gat), .A2(G233gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n237), .A2(new_n239), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n237), .A2(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(new_n234), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n240), .ZN(new_n246));
  XOR2_X1   g045(.A(G183gat), .B(G211gat), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n243), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n243), .B2(new_n246), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n233), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n243), .A2(new_n246), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n243), .A2(new_n246), .A3(new_n248), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n232), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G43gat), .B(G50gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT15), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT89), .B(G29gat), .Z(new_n261));
  INV_X1    g060(.A(G29gat), .ZN(new_n262));
  INV_X1    g061(.A(G36gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT14), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT14), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n265), .B1(G29gat), .B2(G36gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT91), .ZN(new_n268));
  AOI22_X1  g067(.A1(G36gat), .A2(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n260), .B(new_n269), .C1(new_n268), .C2(new_n267), .ZN(new_n270));
  AOI22_X1  g069(.A1(G36gat), .A2(new_n261), .B1(new_n267), .B2(KEYINPUT88), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(KEYINPUT88), .B2(new_n267), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT15), .A3(new_n257), .ZN(new_n273));
  AND2_X1   g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n210), .A2(new_n207), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G229gat), .A2(G233gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT13), .Z(new_n278));
  AND3_X1   g077(.A1(new_n276), .A2(KEYINPUT95), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT95), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(KEYINPUT17), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n282), .B(new_n275), .C1(new_n274), .C2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n274), .A2(new_n275), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(KEYINPUT18), .A3(new_n277), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n284), .A2(new_n277), .A3(new_n285), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT18), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n281), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G113gat), .B(G141gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(G197gat), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT11), .B(G169gat), .Z(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n295), .B(KEYINPUT12), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n281), .A2(new_n298), .A3(new_n287), .A4(new_n290), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G85gat), .A2(G92gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g102(.A1(G99gat), .A2(G106gat), .ZN(new_n304));
  INV_X1    g103(.A(G85gat), .ZN(new_n305));
  INV_X1    g104(.A(G92gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(KEYINPUT8), .A2(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G99gat), .B(G106gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n301), .B1(new_n274), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT102), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n282), .B(new_n311), .C1(new_n274), .C2(new_n283), .ZN(new_n315));
  XOR2_X1   g114(.A(G190gat), .B(G218gat), .Z(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT103), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n321), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT104), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n323), .B2(new_n324), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT106), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n303), .A2(new_n309), .A3(new_n307), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT105), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n222), .A2(new_n228), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n310), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n222), .A2(new_n228), .A3(new_n311), .A4(new_n336), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT10), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n310), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n333), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n339), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n342), .B1(new_n343), .B2(new_n333), .ZN(new_n344));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n344), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n256), .A2(new_n300), .A3(new_n331), .A4(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G227gat), .ZN(new_n353));
  INV_X1    g152(.A(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G183gat), .ZN(new_n357));
  AOI21_X1  g156(.A(G190gat), .B1(new_n357), .B2(KEYINPUT27), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT27), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G183gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(KEYINPUT28), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n361), .B(KEYINPUT72), .Z(new_n362));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n357), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT70), .B(G183gat), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n365), .A2(KEYINPUT71), .A3(new_n369), .A4(new_n358), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n358), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(KEYINPUT27), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n357), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n376), .B2(KEYINPUT70), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT71), .B1(new_n377), .B2(new_n365), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n362), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(KEYINPUT26), .ZN(new_n382));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n383), .B1(new_n380), .B2(KEYINPUT23), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n390), .A2(G169gat), .A3(G176gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G169gat), .ZN(new_n393));
  INV_X1    g192(.A(G176gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT23), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n390), .B1(G169gat), .B2(G176gat), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT65), .A4(new_n383), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT64), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT24), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G190gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n357), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n399), .A2(new_n401), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n397), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n402), .A2(new_n411), .A3(new_n403), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n398), .B1(G183gat), .B2(G190gat), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n411), .B1(new_n402), .B2(new_n403), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT25), .A4(new_n383), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n416), .A2(KEYINPUT67), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT66), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n412), .A3(new_n406), .A4(new_n398), .ZN(new_n421));
  INV_X1    g220(.A(new_n417), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n410), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT68), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT67), .B1(new_n416), .B2(new_n417), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n422), .A3(new_n419), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n410), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n387), .A2(new_n425), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G134gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G127gat), .ZN(new_n433));
  INV_X1    g232(.A(G127gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G134gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G113gat), .B(G120gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(KEYINPUT1), .ZN(new_n438));
  INV_X1    g237(.A(G120gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G113gat), .ZN(new_n440));
  INV_X1    g239(.A(G113gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G120gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G127gat), .B(G134gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n438), .A2(new_n446), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n387), .A2(new_n425), .A3(new_n449), .A4(new_n430), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n356), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(G71gat), .B(G99gat), .Z(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G43gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT33), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n428), .A2(new_n429), .A3(new_n410), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n429), .B1(new_n428), .B2(new_n410), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n449), .B1(new_n463), .B2(new_n387), .ZN(new_n464));
  INV_X1    g263(.A(new_n450), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n355), .B(new_n456), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n466), .B2(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n460), .B1(new_n467), .B2(new_n453), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT74), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT73), .B(new_n456), .C1(new_n451), .C2(KEYINPUT33), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n451), .A2(new_n452), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n460), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n448), .A2(new_n356), .A3(new_n450), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT34), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT34), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n448), .A2(new_n477), .A3(new_n356), .A4(new_n450), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT75), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n469), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n479), .B1(new_n472), .B2(new_n460), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n487));
  INV_X1    g286(.A(new_n479), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n460), .B(new_n479), .C1(new_n467), .C2(new_n453), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  AOI211_X1 g291(.A(KEYINPUT76), .B(KEYINPUT36), .C1(new_n489), .C2(new_n490), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n486), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G1gat), .B(G29gat), .Z(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G57gat), .B(G85gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n501));
  OR2_X1    g300(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(G141gat), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G148gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(G141gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G155gat), .A2(G162gat), .ZN(new_n509));
  INV_X1    g308(.A(G155gat), .ZN(new_n510));
  INV_X1    g309(.A(G162gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n509), .B1(new_n512), .B2(KEYINPUT2), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT2), .ZN(new_n514));
  INV_X1    g313(.A(G141gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G148gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n506), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n512), .A2(new_n509), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n508), .A2(new_n513), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n449), .B1(new_n501), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n521), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n513), .B1(new_n523), .B2(new_n506), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT79), .B1(new_n526), .B2(KEYINPUT3), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n528));
  AOI211_X1 g327(.A(new_n528), .B(new_n501), .C1(new_n524), .C2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n520), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n526), .A2(new_n531), .A3(new_n447), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT4), .B1(new_n449), .B2(new_n519), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G225gat), .A2(G233gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT80), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT5), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n526), .B(new_n447), .ZN(new_n539));
  INV_X1    g338(.A(new_n535), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n530), .A2(new_n534), .A3(new_n538), .A4(new_n535), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n537), .B1(new_n536), .B2(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n500), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n536), .A2(new_n541), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT80), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(new_n499), .A3(new_n543), .A4(new_n542), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT82), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT82), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n546), .A2(new_n550), .A3(new_n553), .A4(new_n547), .ZN(new_n554));
  OAI211_X1 g353(.A(KEYINPUT6), .B(new_n500), .C1(new_n544), .C2(new_n545), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G8gat), .B(G36gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT22), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n561), .A2(KEYINPUT77), .B1(G211gat), .B2(G218gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(KEYINPUT77), .B2(new_n561), .ZN(new_n563));
  XNOR2_X1  g362(.A(G197gat), .B(G204gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G211gat), .B(G218gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  AOI22_X1  g366(.A1(new_n426), .A2(new_n427), .B1(new_n409), .B2(new_n408), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n568), .B1(new_n379), .B2(new_n386), .ZN(new_n569));
  AND2_X1   g368(.A1(G226gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT29), .ZN(new_n571));
  AOI221_X4 g370(.A(new_n567), .B1(new_n569), .B2(new_n570), .C1(new_n431), .C2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n565), .B(new_n566), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n377), .A2(new_n365), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n371), .A3(new_n370), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n385), .B1(new_n577), .B2(new_n362), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n571), .B1(new_n578), .B2(new_n568), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n387), .A2(new_n425), .A3(new_n430), .A4(new_n570), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n573), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n560), .B1(new_n572), .B2(new_n581), .ZN(new_n582));
  AND4_X1   g381(.A1(new_n387), .A2(new_n425), .A3(new_n430), .A4(new_n570), .ZN(new_n583));
  INV_X1    g382(.A(new_n571), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n567), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n425), .A2(new_n430), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n571), .B1(new_n587), .B2(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n570), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n573), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n590), .A3(new_n559), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(KEYINPUT30), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n572), .A2(new_n581), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT30), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n559), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n556), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G78gat), .B(G106gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT31), .B(G50gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n573), .A2(KEYINPUT29), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n526), .B1(new_n602), .B2(KEYINPUT3), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n524), .A2(new_n501), .A3(new_n525), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT29), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n573), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G22gat), .ZN(new_n609));
  INV_X1    g408(.A(G228gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(new_n354), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n567), .A2(new_n605), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n519), .B1(new_n612), .B2(new_n501), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n613), .B2(KEYINPUT83), .ZN(new_n614));
  INV_X1    g413(.A(G22gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n603), .A2(new_n615), .A3(new_n607), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n609), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n609), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n601), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n614), .ZN(new_n620));
  INV_X1    g419(.A(new_n616), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n615), .B1(new_n603), .B2(new_n607), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n609), .A2(new_n614), .A3(new_n616), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n600), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n619), .A2(new_n625), .A3(KEYINPUT84), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT84), .B1(new_n619), .B2(new_n625), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n597), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT85), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n604), .A2(new_n447), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n528), .B1(new_n519), .B2(new_n501), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n526), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n531), .B1(new_n526), .B2(new_n447), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n449), .A2(new_n519), .A3(KEYINPUT4), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n631), .B(new_n540), .C1(new_n635), .C2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n535), .B1(new_n530), .B2(new_n534), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT39), .B1(new_n539), .B2(new_n540), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n639), .B(new_n499), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n630), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n630), .A3(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n549), .A2(new_n543), .A3(new_n542), .ZN(new_n648));
  INV_X1    g447(.A(new_n642), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n648), .A2(new_n500), .B1(new_n649), .B2(KEYINPUT40), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n592), .A2(new_n595), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n642), .A2(new_n630), .A3(new_n643), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n644), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n649), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n546), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n658), .A2(KEYINPUT86), .A3(new_n595), .A4(new_n592), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n619), .A2(new_n625), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT38), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n573), .B1(new_n583), .B2(new_n585), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n588), .A2(new_n567), .A3(new_n589), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT37), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n559), .B1(new_n586), .B2(new_n590), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT37), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n559), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n663), .B(new_n666), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n670), .A2(new_n551), .A3(new_n555), .A4(new_n591), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n559), .B1(new_n593), .B2(new_n668), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT37), .B1(new_n572), .B2(new_n581), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n663), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n662), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n629), .B1(new_n660), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n494), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n555), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n551), .B2(KEYINPUT82), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n680), .A2(new_n554), .B1(new_n595), .B2(new_n592), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n483), .A2(new_n661), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n482), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT35), .ZN(new_n684));
  INV_X1    g483(.A(new_n490), .ZN(new_n685));
  NOR4_X1   g484(.A1(new_n685), .A2(new_n483), .A3(KEYINPUT35), .A4(new_n661), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n551), .A2(new_n555), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n596), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT87), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT87), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n596), .A2(new_n690), .A3(new_n687), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n686), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n352), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n494), .A2(new_n677), .B1(new_n684), .B2(new_n693), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT107), .B1(new_n698), .B2(new_n351), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n556), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  INV_X1    g503(.A(new_n596), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  NAND3_X1  g505(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n697), .A2(new_n699), .ZN(new_n710));
  OAI21_X1  g509(.A(G8gat), .B1(new_n710), .B2(new_n596), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n707), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n704), .B(new_n709), .C1(new_n712), .C2(new_n708), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n708), .B1(new_n711), .B2(new_n707), .ZN(new_n714));
  INV_X1    g513(.A(new_n709), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT108), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1325gat));
  INV_X1    g516(.A(G15gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n710), .A2(new_n718), .A3(new_n494), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n710), .B2(new_n491), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(KEYINPUT109), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(G1326gat));
  NAND2_X1  g522(.A1(new_n700), .A2(new_n628), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT110), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT43), .B(G22gat), .Z(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1327gat));
  AND2_X1   g526(.A1(new_n251), .A2(new_n255), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n300), .A3(new_n350), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n698), .A2(new_n729), .A3(new_n331), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n556), .A2(new_n261), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n484), .B1(new_n685), .B2(new_n483), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT76), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n491), .A2(new_n487), .A3(new_n484), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n676), .B1(new_n737), .B2(new_n486), .ZN(new_n738));
  AOI22_X1  g537(.A1(KEYINPUT35), .A2(new_n683), .B1(new_n686), .B2(new_n692), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT111), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n735), .A2(new_n736), .B1(new_n482), .B2(new_n485), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n694), .B(new_n741), .C1(new_n742), .C2(new_n676), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n331), .A2(KEYINPUT44), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n698), .B2(new_n331), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n729), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n701), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n261), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n749), .B2(new_n701), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n733), .B1(new_n752), .B2(new_n753), .ZN(G1328gat));
  AOI21_X1  g553(.A(G36gat), .B1(KEYINPUT113), .B2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n730), .A2(new_n705), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n748), .A2(new_n596), .A3(new_n729), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n263), .ZN(G1329gat));
  NAND2_X1  g559(.A1(new_n742), .A2(G43gat), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n748), .A2(new_n729), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n491), .ZN(new_n763));
  AOI21_X1  g562(.A(G43gat), .B1(new_n730), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1330gat));
  INV_X1    g566(.A(G50gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n730), .A2(new_n768), .A3(new_n628), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n748), .A2(new_n662), .A3(new_n729), .ZN(new_n770));
  NAND2_X1  g569(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n771));
  OAI221_X1 g570(.A(new_n769), .B1(KEYINPUT114), .B2(KEYINPUT48), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n749), .A2(new_n628), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G50gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n775), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g575(.A1(new_n740), .A2(new_n743), .ZN(new_n777));
  NOR4_X1   g576(.A1(new_n728), .A2(new_n300), .A3(new_n330), .A4(new_n350), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n556), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT97), .B(G57gat), .Z(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1332gat));
  OAI22_X1  g581(.A1(new_n779), .A2(new_n596), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(KEYINPUT49), .B(G64gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n777), .A2(new_n705), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT115), .Z(G1333gat));
  NAND4_X1  g586(.A1(new_n778), .A2(new_n740), .A3(new_n763), .A4(new_n743), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  AOI21_X1  g588(.A(G71gat), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n494), .A2(new_n217), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n778), .A2(new_n740), .A3(new_n743), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT50), .ZN(G1334gat));
  INV_X1    g595(.A(new_n628), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(new_n218), .ZN(G1335gat));
  INV_X1    g598(.A(new_n300), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n251), .A2(new_n255), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n350), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n747), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n556), .ZN(new_n804));
  INV_X1    g603(.A(new_n801), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n330), .C1(new_n738), .C2(new_n739), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n695), .A2(KEYINPUT51), .A3(new_n330), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n701), .A2(new_n305), .A3(new_n349), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  AOI21_X1  g612(.A(new_n331), .B1(new_n678), .B2(new_n694), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n814), .B2(new_n805), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT118), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n808), .A2(new_n809), .A3(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n350), .A2(G92gat), .A3(new_n596), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n802), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n745), .B2(new_n746), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n306), .B1(new_n822), .B2(new_n705), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825));
  INV_X1    g624(.A(new_n819), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n811), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n824), .B1(new_n827), .B2(new_n823), .ZN(G1337gat));
  OAI21_X1  g627(.A(G99gat), .B1(new_n803), .B2(new_n494), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n350), .A2(new_n491), .A3(G99gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n811), .B2(new_n830), .ZN(G1338gat));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n747), .A2(new_n628), .A3(new_n802), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n350), .A2(G106gat), .A3(new_n662), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n818), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n833), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n836), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n833), .ZN(new_n840));
  INV_X1    g639(.A(G106gat), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n822), .B2(new_n661), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n832), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n816), .A2(new_n818), .A3(new_n836), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n822), .B2(new_n628), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT53), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G106gat), .B1(new_n803), .B2(new_n662), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n810), .B2(new_n836), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n851), .ZN(G1339gat));
  NOR2_X1   g651(.A1(new_n344), .A2(new_n348), .ZN(new_n853));
  XOR2_X1   g652(.A(KEYINPUT120), .B(KEYINPUT54), .Z(new_n854));
  OAI211_X1 g653(.A(new_n333), .B(new_n854), .C1(new_n340), .C2(new_n341), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n348), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n855), .A2(KEYINPUT121), .A3(new_n348), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n340), .A2(new_n341), .A3(new_n333), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n342), .A2(KEYINPUT54), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n858), .A2(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n853), .B1(new_n862), .B2(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n860), .ZN(new_n864));
  INV_X1    g663(.A(new_n859), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT121), .B1(new_n855), .B2(new_n348), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n300), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n286), .A2(new_n277), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n276), .A2(new_n278), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n295), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n299), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n349), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n330), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  AND4_X1   g675(.A1(new_n330), .A2(new_n874), .A3(new_n863), .A4(new_n869), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n330), .A2(new_n874), .A3(new_n863), .A4(new_n869), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n297), .A2(new_n299), .B1(new_n867), .B2(new_n868), .ZN(new_n881));
  AOI22_X1  g680(.A1(new_n881), .A2(new_n863), .B1(new_n349), .B2(new_n874), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n879), .B(new_n880), .C1(new_n882), .C2(new_n330), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n728), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n256), .A2(new_n800), .A3(new_n331), .A4(new_n350), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n482), .A2(new_n682), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(new_n701), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT123), .A3(new_n596), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT123), .B1(new_n888), .B2(new_n596), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n441), .B(new_n300), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n491), .A2(new_n628), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n705), .A2(new_n556), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n800), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(G1340gat));
  OAI211_X1 g696(.A(new_n439), .B(new_n349), .C1(new_n889), .C2(new_n890), .ZN(new_n898));
  OAI21_X1  g697(.A(G120gat), .B1(new_n895), .B2(new_n350), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1341gat));
  OAI21_X1  g699(.A(G127gat), .B1(new_n895), .B2(new_n728), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n888), .A2(new_n434), .A3(new_n596), .A4(new_n256), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1342gat));
  NOR2_X1   g702(.A1(new_n331), .A2(new_n705), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n432), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g705(.A(G134gat), .B1(new_n895), .B2(new_n331), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G1343gat));
  NAND4_X1  g708(.A1(new_n886), .A2(new_n701), .A3(new_n494), .A4(new_n661), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n705), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n515), .A3(new_n300), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n662), .B1(new_n884), .B2(new_n885), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n494), .A2(new_n894), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n728), .B1(new_n876), .B2(new_n877), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n797), .B1(new_n918), .B2(new_n885), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n916), .A2(new_n800), .A3(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n912), .B(new_n913), .C1(new_n921), .C2(new_n515), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n915), .B2(new_n914), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n515), .B1(new_n923), .B2(new_n300), .ZN(new_n924));
  NOR4_X1   g723(.A1(new_n910), .A2(G141gat), .A3(new_n705), .A4(new_n800), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT58), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n922), .A2(new_n926), .ZN(G1344gat));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n916), .A2(new_n350), .A3(new_n920), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n521), .A2(new_n522), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n932), .B1(KEYINPUT57), .B2(new_n919), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n349), .A3(new_n917), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n928), .A2(new_n505), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n911), .A2(new_n930), .A3(new_n349), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n936), .A3(new_n937), .ZN(G1345gat));
  INV_X1    g737(.A(new_n923), .ZN(new_n939));
  OAI21_X1  g738(.A(G155gat), .B1(new_n939), .B2(new_n728), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n510), .A3(new_n256), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(G162gat), .B1(new_n939), .B2(new_n331), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n904), .A2(new_n511), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n910), .B2(new_n944), .ZN(G1347gat));
  AOI21_X1  g744(.A(new_n701), .B1(new_n884), .B2(new_n885), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n887), .A2(new_n705), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT124), .Z(new_n948));
  AND2_X1   g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n393), .A3(new_n300), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n701), .A2(new_n596), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n886), .A2(new_n892), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n300), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT125), .A3(G169gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n953), .B2(G169gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(G1348gat));
  INV_X1    g755(.A(new_n952), .ZN(new_n957));
  OAI21_X1  g756(.A(G176gat), .B1(new_n957), .B2(new_n350), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n949), .A2(new_n394), .A3(new_n349), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1349gat));
  AOI21_X1  g759(.A(new_n357), .B1(new_n952), .B2(new_n256), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT60), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n357), .A2(KEYINPUT27), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n256), .A2(new_n964), .A3(new_n360), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n966), .ZN(new_n968));
  OAI21_X1  g767(.A(KEYINPUT60), .B1(new_n968), .B2(new_n961), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1350gat));
  NAND3_X1  g769(.A1(new_n949), .A2(new_n405), .A3(new_n330), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n952), .A2(new_n330), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(G190gat), .ZN(new_n974));
  AOI211_X1 g773(.A(KEYINPUT61), .B(new_n405), .C1(new_n952), .C2(new_n330), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(G1351gat));
  AND4_X1   g775(.A1(new_n494), .A2(new_n946), .A3(new_n705), .A4(new_n661), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n300), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n494), .A2(new_n951), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n933), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n300), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  OAI21_X1  g782(.A(G204gat), .B1(new_n980), .B2(new_n350), .ZN(new_n984));
  NAND2_X1  g783(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n350), .A2(G204gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n977), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n977), .A2(new_n986), .ZN(new_n988));
  XNOR2_X1  g787(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(G1353gat));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n992), .A3(new_n256), .ZN(new_n993));
  AOI211_X1 g792(.A(new_n915), .B(new_n662), .C1(new_n884), .C2(new_n885), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n919), .A2(KEYINPUT57), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n256), .B(new_n979), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  AOI21_X1  g798(.A(G218gat), .B1(new_n977), .B2(new_n330), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n330), .A2(G218gat), .ZN(new_n1001));
  XOR2_X1   g800(.A(new_n1001), .B(KEYINPUT127), .Z(new_n1002));
  AOI21_X1  g801(.A(new_n1000), .B1(new_n981), .B2(new_n1002), .ZN(G1355gat));
endmodule


