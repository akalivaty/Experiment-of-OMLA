//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G137), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(G131), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n200), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n200), .A2(new_n204), .B1(new_n202), .B2(G128), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n198), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT0), .A4(G128), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT0), .B(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n194), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G116), .B(G119), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT2), .B(G113), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(new_n213), .B2(new_n219), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(G237), .A2(G953), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G210), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT27), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT26), .B(G101), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n239));
  INV_X1    g053(.A(new_n235), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n220), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT30), .B1(new_n213), .B2(new_n219), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n225), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT64), .B1(new_n208), .B2(new_n200), .ZN(new_n245));
  AND4_X1   g059(.A1(KEYINPUT64), .A2(new_n200), .A3(new_n202), .A4(new_n204), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n212), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n198), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n216), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n218), .A2(new_n194), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(new_n224), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n240), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n238), .A2(new_n239), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G902), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n240), .A2(new_n239), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n220), .B2(new_n225), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n228), .B2(new_n259), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n237), .B(new_n258), .C1(new_n261), .C2(new_n236), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G472), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n213), .A2(new_n219), .A3(KEYINPUT30), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n241), .B1(new_n249), .B2(new_n252), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n224), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n235), .A3(new_n226), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT31), .ZN(new_n269));
  INV_X1    g083(.A(new_n229), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n226), .B2(new_n227), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n240), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n267), .A2(new_n274), .A3(new_n235), .A4(new_n226), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n269), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n277));
  NOR2_X1   g091(.A1(G472), .A2(G902), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n264), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n264), .B(new_n283), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT16), .ZN(new_n285));
  INV_X1    g099(.A(G140), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(G125), .ZN(new_n288));
  INV_X1    g102(.A(G125), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G140), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n287), .B1(new_n291), .B2(new_n285), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n201), .ZN(new_n293));
  OAI211_X1 g107(.A(G146), .B(new_n287), .C1(new_n291), .C2(new_n285), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(G128), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n298), .B(new_n299), .C1(G119), .C2(new_n199), .ZN(new_n300));
  XNOR2_X1  g114(.A(G119), .B(G128), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT24), .B(G110), .Z(new_n302));
  AOI22_X1  g116(.A1(new_n300), .A2(G110), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n300), .A2(G110), .B1(new_n301), .B2(new_n302), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n305), .B(new_n294), .C1(G146), .C2(new_n291), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G137), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  INV_X1    g123(.A(G234), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(new_n310), .A3(G953), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n308), .B(new_n311), .Z(new_n312));
  XNOR2_X1  g126(.A(new_n307), .B(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G217), .B1(new_n310), .B2(G902), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n257), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n257), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(KEYINPUT25), .ZN(new_n320));
  INV_X1    g134(.A(new_n315), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(KEYINPUT25), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n282), .A2(new_n284), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n282), .A2(KEYINPUT72), .A3(new_n324), .A4(new_n284), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G469), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  INV_X1    g145(.A(G104), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G107), .ZN(new_n333));
  INV_X1    g147(.A(G107), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT3), .A3(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(G107), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n337), .B1(new_n336), .B2(new_n338), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(KEYINPUT4), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n216), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n334), .A2(KEYINPUT3), .A3(G104), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT3), .B1(new_n334), .B2(G104), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT73), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G101), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n342), .B(new_n338), .C1(new_n345), .C2(new_n346), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n334), .B2(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n334), .A2(G104), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n332), .A2(KEYINPUT74), .A3(G107), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G101), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n351), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n247), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n211), .B1(new_n207), .B2(new_n209), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n358), .A2(new_n351), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT10), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n344), .A2(new_n352), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n251), .B1(new_n365), .B2(KEYINPUT77), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n344), .A2(new_n352), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n364), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT78), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT77), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT78), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n251), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n251), .B(KEYINPUT75), .Z(new_n378));
  NOR2_X1   g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  INV_X1    g195(.A(G953), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n382), .A2(G227), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n381), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n359), .A2(new_n247), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n362), .A2(new_n363), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n387), .A2(new_n388), .B1(new_n194), .B2(new_n218), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(KEYINPUT76), .B2(KEYINPUT12), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT76), .B(KEYINPUT12), .Z(new_n391));
  OAI21_X1  g205(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n384), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n330), .B1(new_n395), .B2(new_n257), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT79), .B(G469), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n385), .B1(new_n377), .B2(new_n380), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n380), .A2(new_n392), .A3(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n257), .B(new_n397), .C1(new_n398), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n379), .B1(new_n370), .B2(new_n376), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n399), .B1(new_n403), .B2(new_n385), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT80), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n405), .A3(new_n257), .A4(new_n397), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n396), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT9), .B(G234), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n309), .B1(new_n409), .B2(new_n257), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(G952), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n412), .A2(KEYINPUT87), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n382), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(G234), .B2(G237), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n257), .B1(G234), .B2(G237), .ZN(new_n417));
  INV_X1    g231(.A(G898), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n382), .B1(KEYINPUT21), .B2(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n418), .A2(KEYINPUT21), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n416), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n223), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n221), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n221), .A2(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n297), .A2(G116), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n427), .B(G113), .C1(KEYINPUT5), .C2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n359), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n341), .B2(G101), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n348), .A2(new_n349), .A3(new_n343), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n224), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n436), .B(new_n430), .C1(new_n432), .C2(new_n434), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n250), .A2(G125), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n441), .B1(G125), .B2(new_n362), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT81), .B(G224), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT82), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n442), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n447), .A3(new_n437), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n436), .B(KEYINPUT8), .Z(new_n451));
  NAND2_X1  g265(.A1(new_n429), .A2(new_n426), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n363), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n453), .B2(new_n430), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n444), .A2(KEYINPUT7), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n442), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n442), .A2(new_n455), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n458), .B2(new_n439), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n449), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n450), .B1(new_n449), .B2(new_n459), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n411), .B(new_n424), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G475), .ZN(new_n463));
  XNOR2_X1  g277(.A(G113), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n332), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n291), .B(G146), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n231), .A2(G143), .A3(G214), .ZN(new_n467));
  AOI21_X1  g281(.A(G143), .B1(new_n231), .B2(G214), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT18), .B(G131), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n231), .A2(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n203), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n231), .A2(G143), .A3(G214), .ZN(new_n472));
  NAND2_X1  g286(.A1(KEYINPUT18), .A2(G131), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n466), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(KEYINPUT17), .B(G131), .C1(new_n467), .C2(new_n468), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n293), .A2(new_n476), .A3(new_n294), .ZN(new_n477));
  OAI21_X1  g291(.A(G131), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n192), .A3(new_n472), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n465), .B(new_n475), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(new_n293), .A3(new_n294), .A4(new_n476), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n465), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n257), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n463), .B1(new_n487), .B2(KEYINPUT83), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n475), .B1(new_n477), .B2(new_n481), .ZN(new_n489));
  INV_X1    g303(.A(new_n465), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n491), .B2(new_n482), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n479), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT19), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT19), .B1(new_n288), .B2(new_n290), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n201), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n498), .A3(new_n294), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n465), .B1(new_n499), .B2(new_n475), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n466), .A2(new_n469), .A3(new_n474), .ZN(new_n501));
  INV_X1    g315(.A(new_n477), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n484), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n500), .B1(new_n503), .B2(new_n465), .ZN(new_n504));
  NOR2_X1   g318(.A1(G475), .A2(G902), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT20), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n500), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n482), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT20), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n505), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n488), .A2(new_n494), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G478), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n203), .A2(G128), .ZN(new_n516));
  OAI21_X1  g330(.A(G134), .B1(new_n516), .B2(KEYINPUT13), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n203), .A2(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n199), .A2(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT13), .A4(G134), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G122), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT84), .B1(new_n524), .B2(G116), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n526));
  INV_X1    g340(.A(G116), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(G122), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n525), .A2(new_n528), .B1(G116), .B2(new_n524), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n334), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(G116), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n531), .A2(new_n334), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n523), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT85), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT85), .B1(new_n518), .B2(new_n519), .ZN(new_n537));
  OAI21_X1  g351(.A(G134), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n520), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n535), .A3(new_n188), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n334), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n531), .A2(KEYINPUT14), .B1(G116), .B2(new_n524), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n525), .A2(new_n528), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n334), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n534), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n409), .A2(G217), .A3(new_n382), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n534), .B(new_n551), .C1(new_n543), .C2(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT86), .B(G902), .C1(new_n550), .C2(new_n552), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n515), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n514), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n512), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NOR4_X1   g374(.A1(new_n407), .A2(new_n410), .A3(new_n462), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n329), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT88), .B(G101), .Z(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(G3));
  NAND2_X1  g378(.A1(new_n402), .A2(new_n406), .ZN(new_n565));
  INV_X1    g379(.A(new_n396), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n410), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n462), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n553), .A2(G478), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT33), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT89), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n531), .A2(KEYINPUT14), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n532), .A3(new_n546), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G107), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(new_n542), .A3(new_n541), .A4(new_n538), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n551), .B1(new_n581), .B2(new_n534), .ZN(new_n582));
  INV_X1    g396(.A(new_n552), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n574), .B(new_n577), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n550), .A2(KEYINPUT89), .A3(new_n575), .A4(new_n552), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n513), .A2(G902), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n571), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n512), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT90), .B1(new_n570), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT90), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n462), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n276), .A2(new_n278), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n276), .A2(new_n257), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n324), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n569), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT91), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT34), .B(G104), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NOR3_X1   g416(.A1(new_n407), .A2(new_n598), .A3(new_n410), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n557), .A2(new_n559), .B1(new_n494), .B2(new_n488), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n511), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n510), .B1(new_n509), .B2(new_n505), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT20), .B(new_n506), .C1(new_n508), .C2(new_n482), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n609), .B2(new_n605), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n604), .A2(new_n424), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n612));
  INV_X1    g426(.A(new_n411), .ZN(new_n613));
  INV_X1    g427(.A(new_n461), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n449), .A2(new_n450), .A3(new_n459), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n604), .A2(new_n617), .A3(new_n424), .A4(new_n610), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n612), .A2(KEYINPUT94), .A3(new_n616), .A4(new_n618), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n603), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n334), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n597), .A2(new_n595), .ZN(new_n628));
  INV_X1    g442(.A(new_n312), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n307), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n317), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n320), .B2(new_n322), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n561), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  NOR2_X1   g452(.A1(new_n407), .A2(new_n410), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n282), .A2(new_n284), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n416), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n382), .A2(G900), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n417), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT96), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n644), .A2(KEYINPUT96), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n604), .A2(new_n610), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n616), .A2(new_n633), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n639), .A2(new_n641), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT97), .B(G128), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G30));
  XNOR2_X1  g467(.A(new_n647), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n639), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n614), .A2(new_n615), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n512), .B1(new_n557), .B2(new_n559), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n411), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n228), .A2(new_n259), .ZN(new_n661));
  INV_X1    g475(.A(new_n260), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n257), .B1(new_n663), .B2(new_n235), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n267), .A2(new_n226), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n235), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT98), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n280), .B2(new_n279), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n634), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n660), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n656), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NOR4_X1   g491(.A1(new_n407), .A2(new_n640), .A3(new_n410), .A4(new_n649), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n589), .A2(new_n647), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n639), .A2(new_n641), .A3(new_n650), .A4(new_n681), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NOR2_X1   g500(.A1(new_n594), .A2(new_n325), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n404), .A2(new_n257), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n565), .A2(new_n568), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n402), .A2(new_n406), .B1(G469), .B2(new_n688), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(KEYINPUT101), .A3(new_n568), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n687), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n687), .A2(new_n692), .A3(KEYINPUT102), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  AND2_X1   g515(.A1(new_n692), .A2(new_n694), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n325), .B1(new_n621), .B2(new_n622), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT103), .B(G116), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G18));
  AND4_X1   g520(.A1(new_n568), .A2(new_n565), .A3(new_n616), .A4(new_n689), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n633), .A2(new_n424), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n640), .A2(new_n560), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NAND2_X1  g525(.A1(new_n663), .A2(KEYINPUT28), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n235), .B1(new_n712), .B2(new_n237), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n269), .A2(new_n275), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n278), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n323), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n597), .A2(KEYINPUT104), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n597), .A2(KEYINPUT104), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n616), .A2(new_n659), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n423), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n702), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  OAI211_X1 g537(.A(new_n715), .B(new_n633), .C1(new_n717), .C2(new_n718), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n680), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n693), .A3(new_n568), .A4(new_n616), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT105), .B(G125), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G27));
  NAND2_X1  g542(.A1(new_n281), .A2(new_n716), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT108), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n730), .A2(new_n731), .A3(new_n680), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n657), .A2(new_n613), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n568), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n567), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n407), .B2(new_n735), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n732), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n325), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n733), .B1(new_n567), .B2(new_n736), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n407), .A2(new_n735), .A3(KEYINPUT106), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n741), .B(new_n681), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n731), .B1(new_n744), .B2(KEYINPUT107), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n325), .B1(new_n737), .B2(new_n738), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n746), .B1(new_n747), .B2(new_n681), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  OAI211_X1 g564(.A(new_n741), .B(new_n648), .C1(new_n742), .C2(new_n743), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n395), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n386), .A2(KEYINPUT45), .A3(new_n394), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n565), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n568), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(G475), .B1(new_n492), .B2(new_n493), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n766));
  OAI22_X1  g580(.A1(new_n765), .A2(new_n766), .B1(new_n607), .B2(new_n608), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n588), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(KEYINPUT109), .B2(KEYINPUT43), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n628), .A3(new_n633), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT110), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n734), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT110), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n764), .A2(new_n654), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(new_n734), .ZN(new_n780));
  NOR4_X1   g594(.A1(new_n641), .A2(new_n324), .A3(new_n680), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n763), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n763), .A2(new_n782), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(new_n740), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n325), .B(new_n680), .C1(new_n737), .C2(new_n738), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT42), .B1(new_n789), .B2(new_n746), .ZN(new_n790));
  INV_X1    g604(.A(new_n748), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n257), .B1(new_n582), .B2(new_n583), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT86), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n514), .B1(new_n794), .B2(new_n558), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n556), .A2(new_n515), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n557), .A2(new_n798), .A3(new_n559), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT114), .B1(new_n800), .B2(new_n512), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n802), .B(new_n767), .C1(new_n797), .C2(new_n799), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n570), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n512), .B2(new_n588), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n573), .B(new_n576), .C1(new_n550), .C2(new_n552), .ZN(new_n809));
  INV_X1    g623(.A(new_n585), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n587), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n571), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n767), .A3(KEYINPUT111), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n806), .B1(new_n570), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n808), .A2(new_n814), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n462), .A3(KEYINPUT112), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n820), .B(new_n570), .C1(new_n801), .C2(new_n803), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n805), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n822), .A2(new_n603), .B1(new_n707), .B2(new_n709), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n692), .B(new_n694), .C1(new_n703), .C2(new_n721), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n561), .B1(new_n329), .B2(new_n635), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n488), .A2(new_n494), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n633), .A2(new_n827), .A3(new_n610), .A4(new_n647), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n780), .A2(new_n800), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n639), .A2(new_n829), .A3(new_n641), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n725), .B1(new_n742), .B2(new_n743), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n751), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n832), .A3(new_n699), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n792), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n697), .B2(new_n698), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n749), .A3(new_n837), .A4(new_n832), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n651), .A2(new_n726), .ZN(new_n840));
  INV_X1    g654(.A(new_n647), .ZN(new_n841));
  OR4_X1    g655(.A1(new_n569), .A2(new_n841), .A3(new_n671), .A4(new_n720), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n679), .B1(new_n678), .B2(new_n681), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n840), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n651), .A2(new_n726), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n682), .B2(new_n684), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n842), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n840), .A2(new_n849), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n851), .B(new_n855), .C1(new_n834), .C2(new_n838), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n792), .A2(new_n833), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n852), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n851), .B1(new_n834), .B2(new_n838), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(KEYINPUT53), .ZN(new_n864));
  INV_X1    g678(.A(new_n719), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n771), .A2(new_n416), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n690), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n658), .A2(new_n411), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n324), .A2(new_n416), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n690), .A2(new_n670), .A3(new_n780), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n813), .A2(new_n767), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n873), .A2(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n869), .A2(new_n734), .A3(new_n866), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n565), .A2(new_n689), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n568), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n785), .A2(new_n784), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n868), .A2(new_n734), .ZN(new_n885));
  OAI221_X1 g699(.A(new_n878), .B1(new_n724), .B2(new_n881), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n881), .A2(new_n730), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n890), .A2(KEYINPUT118), .A3(KEYINPUT48), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n876), .A2(new_n589), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n415), .B1(new_n868), .B2(new_n707), .ZN(new_n893));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n892), .B(new_n893), .C1(new_n890), .C2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n888), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n857), .A2(new_n864), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n412), .A2(new_n382), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n901));
  INV_X1    g715(.A(new_n768), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n716), .A2(new_n568), .A3(new_n411), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n670), .A2(new_n658), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n900), .A2(KEYINPUT119), .A3(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(G75));
  NAND2_X1  g725(.A1(new_n440), .A2(new_n448), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(new_n446), .Z(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n861), .B1(new_n863), .B2(KEYINPUT53), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n915), .A2(G210), .A3(G902), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n916), .B2(KEYINPUT56), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n382), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n915), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT120), .B1(new_n921), .B2(new_n257), .ZN(new_n922));
  INV_X1    g736(.A(new_n450), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n915), .A2(new_n924), .A3(G902), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n927));
  NOR2_X1   g741(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n926), .B2(new_n928), .ZN(G51));
  XOR2_X1   g743(.A(new_n757), .B(KEYINPUT57), .Z(new_n930));
  NOR2_X1   g744(.A1(new_n921), .A2(new_n862), .ZN(new_n931));
  INV_X1    g745(.A(new_n864), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n404), .ZN(new_n934));
  INV_X1    g748(.A(new_n756), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n922), .A2(new_n935), .A3(new_n925), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n918), .B1(new_n934), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT122), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n922), .A2(new_n925), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n504), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n922), .A2(new_n509), .A3(new_n925), .A4(new_n939), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n941), .A2(new_n919), .A3(new_n942), .ZN(G60));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n857), .B2(new_n864), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(new_n586), .ZN(new_n947));
  INV_X1    g761(.A(new_n945), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n586), .B(new_n948), .C1(new_n931), .C2(new_n932), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n947), .A2(new_n919), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  NAND2_X1  g766(.A1(new_n915), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n313), .B(KEYINPUT123), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n631), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n955), .B(new_n919), .C1(new_n956), .C2(new_n953), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G66));
  NAND2_X1  g773(.A1(new_n443), .A2(G953), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n421), .B(new_n960), .C1(new_n836), .C2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n912), .B1(G898), .B2(new_n382), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  NAND2_X1  g777(.A1(new_n786), .A2(new_n778), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n730), .A2(new_n720), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n764), .A2(new_n654), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n848), .A2(new_n966), .A3(new_n751), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n749), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n643), .B1(new_n969), .B2(new_n382), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n265), .A2(new_n266), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n496), .A2(new_n497), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n382), .B1(G227), .B2(G900), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  OAI22_X1  g789(.A1(new_n970), .A2(new_n973), .B1(KEYINPUT125), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n329), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n801), .A2(new_n803), .A3(new_n815), .ZN(new_n978));
  NOR4_X1   g792(.A1(new_n977), .A2(new_n655), .A3(new_n780), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n964), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n676), .A2(new_n848), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n980), .A2(new_n982), .A3(KEYINPUT124), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n382), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n976), .B1(new_n989), .B2(new_n973), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n975), .A2(KEYINPUT125), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(G72));
  NAND3_X1  g806(.A1(new_n986), .A2(new_n836), .A3(new_n987), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n667), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n255), .A2(new_n268), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n996), .B(new_n999), .C1(new_n853), .C2(new_n856), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n968), .A2(new_n749), .A3(new_n836), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n996), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n665), .A2(new_n235), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n918), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n998), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT127), .ZN(G57));
endmodule


