//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n461), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n464), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n468), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(new_n467), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n461), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n481), .A2(KEYINPUT68), .A3(G124), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n481), .B2(G124), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n473), .B1(new_n474), .B2(new_n475), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(G162));
  NAND2_X1  g060(.A1(new_n481), .A2(G126), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n490), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n461), .B2(G114), .ZN(new_n496));
  AND4_X1   g071(.A1(new_n487), .A2(new_n494), .A3(new_n492), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n486), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(new_n479), .A3(G138), .A4(new_n461), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n466), .A2(KEYINPUT4), .A3(G138), .A4(new_n461), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT72), .Z(new_n511));
  INV_X1    g086(.A(new_n507), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n511), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(new_n509), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT5), .B(G543), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  NAND2_X1  g104(.A1(new_n509), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n514), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n517), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  AOI22_X1  g111(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n517), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT73), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n525), .A2(new_n507), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G81), .B1(new_n509), .B2(G43), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n509), .A2(G53), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT9), .Z(new_n551));
  INV_X1    g126(.A(G91), .ZN(new_n552));
  XNOR2_X1  g127(.A(KEYINPUT75), .B(G65), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n513), .A2(new_n553), .B1(G78), .B2(G543), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n514), .A2(new_n552), .B1(new_n554), .B2(new_n517), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  OR2_X1    g133(.A1(new_n511), .A2(new_n518), .ZN(G303));
  NAND2_X1  g134(.A1(new_n540), .A2(G87), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n509), .A2(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(G288));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n525), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n540), .A2(G86), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n509), .A2(G48), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n571), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n509), .A2(G47), .ZN(new_n575));
  INV_X1    g150(.A(G85), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n514), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n517), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n540), .A2(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  NAND2_X1  g159(.A1(new_n513), .A2(G66), .ZN(new_n585));
  INV_X1    g160(.A(G79), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT77), .B1(new_n586), .B2(new_n508), .ZN(new_n587));
  OR3_X1    g162(.A1(new_n586), .A2(new_n508), .A3(KEYINPUT77), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n509), .B2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n582), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n556), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(new_n556), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n592), .B1(new_n598), .B2(G860), .ZN(G148));
  NAND2_X1  g174(.A1(new_n592), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(KEYINPUT78), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(KEYINPUT78), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n602), .B(new_n603), .C1(G868), .C2(new_n542), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n472), .A2(G2104), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(G2100), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n472), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n481), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n461), .A2(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT79), .B(G2096), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n610), .A2(new_n611), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(G2443), .B(G2446), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT80), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT18), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(new_n609), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1991), .B(G1996), .Z(new_n649));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT19), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  MUX2_X1   g235(.A(new_n660), .B(new_n659), .S(new_n652), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT83), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n649), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  INV_X1    g247(.A(new_n667), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n649), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n675), .A3(new_n668), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n671), .A2(new_n676), .A3(new_n678), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(G229));
  NAND2_X1  g257(.A1(new_n481), .A2(G129), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n689));
  INV_X1    g264(.A(G141), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n688), .B(new_n689), .C1(new_n467), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(G32), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT27), .B(G1996), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G20), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT23), .Z(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G299), .B2(G16), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1956), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G19), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n539), .A2(new_n541), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G1341), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(G1341), .ZN(new_n710));
  AND4_X1   g285(.A1(new_n698), .A2(new_n703), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n693), .A2(G33), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n461), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n714), .B(new_n716), .C1(G139), .C2(new_n472), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n717), .B2(new_n693), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G2072), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n592), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G4), .B2(G16), .ZN(new_n722));
  INV_X1    g297(.A(G1348), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n481), .A2(G128), .ZN(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n728));
  INV_X1    g303(.A(G140), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n728), .C1(new_n729), .C2(new_n467), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n693), .A2(G26), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT31), .B(G11), .Z(new_n737));
  INV_X1    g312(.A(G28), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT30), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT90), .Z(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n738), .B2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n742), .B1(new_n693), .B2(new_n616), .C1(new_n695), .C2(new_n696), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n699), .A2(G5), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G301), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  NOR2_X1   g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n693), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT87), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G160), .B2(G29), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2084), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n699), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n699), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G1966), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(G2084), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n747), .A2(new_n753), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n693), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n693), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n745), .A2(new_n746), .B1(G1966), .B2(new_n755), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n743), .A2(new_n758), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  AND4_X1   g338(.A1(new_n711), .A2(new_n724), .A3(new_n736), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G162), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n693), .A2(G35), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT29), .ZN(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n766), .A2(new_n772), .A3(new_n768), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n770), .A2(new_n771), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n770), .A2(new_n773), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G2090), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n764), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n699), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(G288), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n699), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT33), .B(G1976), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n699), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n699), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G6), .A2(G16), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n572), .A2(new_n573), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT85), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT86), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n788), .A2(new_n789), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n796), .A2(new_n799), .A3(new_n800), .A4(new_n783), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n798), .A2(KEYINPUT34), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n693), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n472), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G119), .ZN(new_n808));
  OR2_X1    g383(.A1(G95), .A2(G2105), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n812), .B2(new_n693), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n699), .A2(G24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n580), .B2(new_n699), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n804), .A2(new_n805), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n804), .A2(new_n822), .A3(new_n805), .A4(new_n819), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n778), .B1(new_n821), .B2(new_n823), .ZN(G311));
  INV_X1    g399(.A(KEYINPUT93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n823), .ZN(new_n826));
  INV_X1    g401(.A(new_n778), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g403(.A(KEYINPUT93), .B(new_n778), .C1(new_n821), .C2(new_n823), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(G150));
  NAND2_X1  g405(.A1(new_n592), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n509), .A2(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n514), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n517), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n542), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n706), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n832), .B(new_n842), .Z(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT39), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT94), .B(G860), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n838), .A2(new_n846), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n730), .B(KEYINPUT96), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n717), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n472), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n481), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n461), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n607), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n854), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G126), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n480), .A2(new_n862), .A3(new_n461), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n494), .A2(new_n492), .A3(new_n496), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT71), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n494), .A2(new_n496), .A3(new_n487), .A4(new_n492), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT95), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT95), .B1(new_n501), .B2(new_n502), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n692), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n812), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n860), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n854), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n616), .B(G160), .ZN(new_n879));
  XNOR2_X1  g454(.A(G162), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n852), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g457(.A(KEYINPUT97), .B(new_n880), .C1(new_n873), .C2(new_n877), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n878), .B2(new_n881), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n851), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n873), .A2(new_n877), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT97), .B1(new_n888), .B2(new_n880), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n878), .A2(new_n852), .A3(new_n881), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n886), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT98), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n887), .A2(new_n893), .A3(KEYINPUT40), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT40), .B1(new_n887), .B2(new_n893), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(G395));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n591), .A2(new_n556), .A3(KEYINPUT99), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n591), .A2(new_n556), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n584), .B(new_n590), .C1(new_n551), .C2(new_n555), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(KEYINPUT99), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n900), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  AOI211_X1 g480(.A(KEYINPUT101), .B(KEYINPUT41), .C1(new_n899), .C2(new_n900), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n902), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n901), .A2(KEYINPUT100), .A3(new_n898), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT100), .B1(new_n898), .B2(new_n901), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n842), .B(new_n600), .ZN(new_n911));
  MUX2_X1   g486(.A(new_n907), .B(new_n910), .S(new_n911), .Z(new_n912));
  NAND2_X1  g487(.A1(G305), .A2(G288), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n792), .A2(new_n780), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G303), .A2(new_n580), .ZN(new_n916));
  NAND2_X1  g491(.A1(G166), .A2(G290), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n916), .A4(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(KEYINPUT102), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n922), .B1(new_n926), .B2(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n912), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(G868), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n929), .B1(G868), .B2(new_n838), .ZN(G295));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n838), .ZN(G331));
  XNOR2_X1  g506(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n898), .A2(new_n901), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n839), .A2(G301), .A3(new_n841), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G301), .B1(new_n839), .B2(new_n841), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(G286), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n842), .A2(G171), .ZN(new_n940));
  AOI21_X1  g515(.A(G168), .B1(new_n940), .B2(new_n936), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(G286), .B1(new_n937), .B2(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(G168), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n942), .B(KEYINPUT104), .C1(new_n907), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n947), .A3(new_n935), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n926), .ZN(new_n950));
  AOI21_X1  g525(.A(G37), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n925), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT102), .B1(new_n919), .B2(new_n920), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n924), .A2(new_n955), .A3(new_n925), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n946), .A2(new_n948), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n933), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n926), .B1(new_n946), .B2(new_n948), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n939), .A2(new_n941), .B1(new_n908), .B2(new_n909), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n935), .A2(new_n897), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n900), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n944), .A3(new_n943), .A4(new_n962), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n954), .A2(new_n956), .A3(new_n960), .A4(new_n963), .ZN(new_n964));
  NOR4_X1   g539(.A1(new_n959), .A2(new_n964), .A3(KEYINPUT43), .A4(G37), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n932), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n951), .A2(new_n957), .A3(new_n933), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n959), .A2(new_n964), .A3(G37), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n967), .B(KEYINPUT44), .C1(new_n933), .C2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G40), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n468), .A2(new_n470), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n501), .A2(new_n502), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n867), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT95), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n503), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT95), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n981), .B2(new_n867), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT45), .ZN(new_n984));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n977), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G2078), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT53), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n870), .A2(new_n992), .A3(new_n985), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n972), .B1(new_n974), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT116), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n870), .A2(new_n992), .A3(new_n985), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n498), .B2(new_n503), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n972), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n746), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n870), .B2(new_n985), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n985), .B(new_n976), .C1(new_n498), .C2(new_n503), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n972), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT53), .A3(new_n989), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1001), .A2(KEYINPUT123), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT123), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n991), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G171), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G288), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT52), .B1(G288), .B2(new_n1011), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n870), .A2(new_n972), .A3(new_n985), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1015), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT110), .B1(new_n1015), .B2(G8), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1013), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n570), .A2(G1981), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(G1981), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT49), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1015), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1015), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1012), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1018), .B(new_n1025), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(G166), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(G160), .A2(G40), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1040), .B1(new_n992), .B2(new_n974), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n870), .A2(new_n985), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT50), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1041), .A2(new_n771), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n977), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n983), .B1(new_n982), .B2(KEYINPUT45), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT109), .B(G1971), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1044), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1039), .B1(new_n1051), .B2(new_n1036), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n988), .A2(new_n1049), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n993), .A2(new_n994), .A3(G2090), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1038), .B(G8), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1033), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1010), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n996), .A2(new_n998), .A3(new_n1060), .A4(new_n972), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT121), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT121), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G168), .A2(new_n1036), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1063), .A2(KEYINPUT122), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1059), .A2(new_n1064), .A3(new_n1061), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1064), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1073));
  OAI21_X1  g648(.A(G168), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1036), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1062), .A2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1066), .A2(KEYINPUT51), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1074), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT62), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1081));
  AOI21_X1  g656(.A(G286), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1076), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1057), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1025), .A2(new_n1011), .A3(new_n780), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1088), .A2(new_n1021), .B1(new_n1029), .B2(new_n1028), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1055), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1033), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1093));
  NAND3_X1  g668(.A1(new_n1062), .A2(G8), .A3(G168), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1056), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT113), .ZN(new_n1096));
  OAI21_X1  g671(.A(G8), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1038), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1090), .A2(new_n1032), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1094), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1100), .A2(KEYINPUT63), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1093), .C1(new_n1056), .C2(new_n1094), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n988), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n556), .B(KEYINPUT57), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1110), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT61), .A3(new_n1114), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1996), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n988), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1015), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n706), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT119), .B(new_n706), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1130), .A2(KEYINPUT59), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1122), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n592), .B2(KEYINPUT120), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1015), .A2(G2067), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT115), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n995), .A2(new_n723), .A3(new_n1000), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1138), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n591), .ZN(new_n1147));
  OAI221_X1 g722(.A(new_n1138), .B1(KEYINPUT120), .B2(new_n592), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT117), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1137), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n1148), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n592), .A3(new_n1151), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT118), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1150), .A2(new_n1156), .A3(new_n592), .A4(new_n1151), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1157), .A3(new_n1120), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1136), .A2(new_n1153), .B1(new_n1158), .B2(new_n1114), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n469), .A2(KEYINPUT124), .ZN(new_n1161));
  OAI21_X1  g736(.A(G2105), .B1(new_n469), .B2(KEYINPUT124), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n989), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1163), .A2(new_n468), .A3(new_n1164), .ZN(new_n1165));
  OAI221_X1 g740(.A(new_n1165), .B1(new_n982), .B2(new_n976), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n991), .A2(new_n1001), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1167), .B2(G171), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1001), .A2(KEYINPUT123), .A3(new_n1006), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n990), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1174), .B2(G301), .ZN(new_n1175));
  OAI211_X1 g750(.A(G301), .B(new_n991), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(KEYINPUT125), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1168), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1056), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1174), .A2(G301), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1167), .A2(G171), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1160), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1084), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1092), .B(new_n1106), .C1(new_n1159), .C2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n982), .A2(new_n1040), .A3(new_n976), .ZN(new_n1186));
  INV_X1    g761(.A(G1986), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n580), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g763(.A(new_n1188), .B(KEYINPUT107), .Z(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1190), .B1(new_n1187), .B2(new_n580), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n730), .B(G2067), .Z(new_n1192));
  XNOR2_X1  g767(.A(new_n692), .B(G1996), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n812), .A2(new_n814), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n812), .A2(new_n814), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1186), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1185), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1186), .A2(new_n1123), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT46), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1199), .B(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1192), .A2(new_n692), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1204), .A2(new_n1186), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  XOR2_X1   g781(.A(new_n1206), .B(KEYINPUT47), .Z(new_n1207));
  NAND2_X1  g782(.A1(new_n1189), .A2(new_n1186), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT127), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT48), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g786(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  AOI211_X1 g787(.A(new_n1211), .B(new_n1212), .C1(new_n1186), .C2(new_n1196), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1214));
  OAI22_X1  g789(.A1(new_n1214), .A2(new_n1194), .B1(G2067), .B2(new_n730), .ZN(new_n1215));
  AOI211_X1 g790(.A(new_n1207), .B(new_n1213), .C1(new_n1186), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1198), .A2(new_n1216), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g792(.A1(new_n958), .A2(new_n965), .ZN(new_n1219));
  INV_X1    g793(.A(G319), .ZN(new_n1220));
  NOR2_X1   g794(.A1(G227), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n634), .B2(new_n635), .ZN(new_n1222));
  AOI21_X1  g796(.A(new_n1222), .B1(new_n680), .B2(new_n681), .ZN(new_n1223));
  AOI21_X1  g797(.A(KEYINPUT98), .B1(new_n891), .B2(new_n892), .ZN(new_n1224));
  AOI211_X1 g798(.A(new_n851), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1219), .A2(new_n1226), .ZN(G308));
  OAI221_X1 g801(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .C1(new_n958), .C2(new_n965), .ZN(G225));
endmodule


