

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n567), .A2(n566), .ZN(G164) );
  NAND2_X1 U554 ( .A1(n685), .A2(n783), .ZN(n720) );
  NOR2_X1 U555 ( .A1(G651), .A2(n632), .ZN(n652) );
  NOR2_X1 U556 ( .A1(G543), .A2(G651), .ZN(n647) );
  NOR2_X2 U557 ( .A1(n549), .A2(n548), .ZN(G160) );
  NOR2_X4 U558 ( .A1(n545), .A2(G2105), .ZN(n887) );
  XOR2_X2 U559 ( .A(G2104), .B(KEYINPUT64), .Z(n545) );
  XOR2_X1 U560 ( .A(G651), .B(KEYINPUT66), .Z(n518) );
  NOR2_X1 U561 ( .A1(G299), .A2(n708), .ZN(n704) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n713) );
  BUF_X1 U563 ( .A(n720), .Z(n733) );
  INV_X1 U564 ( .A(KEYINPUT109), .ZN(n740) );
  XOR2_X1 U565 ( .A(KEYINPUT1), .B(n523), .Z(n650) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  OR2_X1 U567 ( .A1(n632), .A2(n518), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n519), .B(KEYINPUT67), .ZN(n646) );
  NAND2_X1 U569 ( .A1(G78), .A2(n646), .ZN(n521) );
  NAND2_X1 U570 ( .A1(G91), .A2(n647), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U572 ( .A(KEYINPUT71), .B(n522), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n652), .A2(G53), .ZN(n525) );
  NOR2_X1 U574 ( .A1(G543), .A2(n518), .ZN(n523) );
  NAND2_X1 U575 ( .A1(G65), .A2(n650), .ZN(n524) );
  AND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(G299) );
  XNOR2_X1 U578 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n539) );
  NAND2_X1 U579 ( .A1(n647), .A2(G89), .ZN(n528) );
  XNOR2_X1 U580 ( .A(n528), .B(KEYINPUT4), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G76), .A2(n646), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n531), .B(KEYINPUT5), .ZN(n537) );
  XNOR2_X1 U584 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G51), .A2(n652), .ZN(n533) );
  NAND2_X1 U586 ( .A1(G63), .A2(n650), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n535), .B(n534), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n539), .B(n538), .ZN(G168) );
  XOR2_X1 U591 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U592 ( .A1(G101), .A2(n887), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n540), .B(KEYINPUT23), .ZN(n541) );
  XNOR2_X1 U594 ( .A(n541), .B(KEYINPUT65), .ZN(n544) );
  NOR2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XOR2_X1 U596 ( .A(KEYINPUT17), .B(n542), .Z(n886) );
  NAND2_X1 U597 ( .A1(G137), .A2(n886), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n549) );
  AND2_X2 U599 ( .A1(n545), .A2(G2105), .ZN(n882) );
  NAND2_X1 U600 ( .A1(G125), .A2(n882), .ZN(n547) );
  AND2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U602 ( .A1(G113), .A2(n883), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U605 ( .A1(G99), .A2(n887), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G111), .A2(n883), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G135), .A2(n886), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n882), .A2(G123), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n557), .B(KEYINPUT80), .ZN(n981) );
  XNOR2_X1 U614 ( .A(n981), .B(G2096), .ZN(n558) );
  OR2_X1 U615 ( .A1(G2100), .A2(n558), .ZN(G156) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  INV_X1 U619 ( .A(KEYINPUT93), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n882), .A2(G126), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n560), .B(n559), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n883), .A2(G114), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT94), .B(n563), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n887), .A2(G102), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n886), .A2(G138), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n832) );
  NAND2_X1 U631 ( .A1(n832), .A2(G567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n571) );
  NAND2_X1 U634 ( .A1(G56), .A2(n650), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G81), .A2(n647), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT12), .B(n572), .Z(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT73), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G68), .A2(n646), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n652), .A2(G43), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n1016) );
  INV_X1 U645 ( .A(G860), .ZN(n603) );
  OR2_X1 U646 ( .A1(n1016), .A2(n603), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G52), .A2(n652), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT70), .B(n581), .Z(n586) );
  NAND2_X1 U649 ( .A1(G77), .A2(n646), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G90), .A2(n647), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT9), .B(n584), .Z(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n650), .A2(G64), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G66), .A2(n650), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G92), .A2(n647), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G79), .A2(n646), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G54), .A2(n652), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n595), .Z(n596) );
  XNOR2_X2 U664 ( .A(KEYINPUT74), .B(n596), .ZN(n1001) );
  INV_X1 U665 ( .A(G868), .ZN(n666) );
  AND2_X1 U666 ( .A1(n1001), .A2(n666), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n666), .A2(G301), .ZN(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(G284) );
  XNOR2_X1 U669 ( .A(KEYINPUT77), .B(G868), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G286), .A2(n599), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT78), .ZN(n602) );
  NOR2_X1 U672 ( .A1(G299), .A2(G868), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n604), .A2(n1001), .ZN(n605) );
  XNOR2_X1 U676 ( .A(n605), .B(KEYINPUT79), .ZN(n606) );
  XOR2_X1 U677 ( .A(KEYINPUT16), .B(n606), .Z(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n1016), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n1001), .A2(G868), .ZN(n607) );
  NOR2_X1 U680 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U682 ( .A1(n650), .A2(G67), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT84), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G55), .A2(n652), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT85), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G93), .A2(n647), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U689 ( .A1(G80), .A2(n646), .ZN(n616) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(n616), .ZN(n617) );
  NOR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n665) );
  XNOR2_X1 U692 ( .A(n1016), .B(KEYINPUT81), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n1001), .A2(G559), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n620), .B(n619), .ZN(n663) );
  XOR2_X1 U695 ( .A(n663), .B(KEYINPUT82), .Z(n621) );
  NOR2_X1 U696 ( .A1(G860), .A2(n621), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n665), .B(n622), .ZN(G145) );
  XOR2_X1 U698 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n624) );
  NAND2_X1 U699 ( .A1(G73), .A2(n646), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n624), .B(n623), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G48), .A2(n652), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G61), .A2(n650), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n647), .A2(G86), .ZN(n627) );
  XOR2_X1 U705 ( .A(KEYINPUT86), .B(n627), .Z(n628) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G87), .A2(n632), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n650), .A2(n635), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n652), .A2(G49), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U714 ( .A1(n646), .A2(G72), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(KEYINPUT68), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G60), .A2(n650), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G47), .A2(n652), .ZN(n641) );
  XNOR2_X1 U719 ( .A(KEYINPUT69), .B(n641), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n647), .A2(G85), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U723 ( .A1(G75), .A2(n646), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G88), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n657) );
  NAND2_X1 U726 ( .A1(G62), .A2(n650), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(KEYINPUT88), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G50), .A2(n652), .ZN(n653) );
  XOR2_X1 U729 ( .A(KEYINPUT89), .B(n653), .Z(n654) );
  NAND2_X1 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(G166) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(G305), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n665), .B(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(G290), .B(G166), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U737 ( .A(n662), .B(G299), .Z(n898) );
  XNOR2_X1 U738 ( .A(n898), .B(n663), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT90), .B(n669), .Z(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n671), .ZN(n673) );
  XOR2_X1 U746 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n672) );
  XNOR2_X1 U747 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U748 ( .A1(G2072), .A2(n674), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U752 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G96), .A2(n677), .ZN(n836) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n836), .ZN(n681) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U756 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(G108), .A2(n679), .ZN(n837) );
  NAND2_X1 U758 ( .A1(G567), .A2(n837), .ZN(n680) );
  NAND2_X1 U759 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U760 ( .A(KEYINPUT92), .B(n682), .Z(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n684) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n835) );
  NAND2_X1 U764 ( .A1(n835), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  INV_X1 U766 ( .A(G301), .ZN(G171) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n782) );
  INV_X1 U768 ( .A(n782), .ZN(n685) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n783) );
  INV_X1 U770 ( .A(G1996), .ZN(n686) );
  NOR2_X1 U771 ( .A1(n720), .A2(n686), .ZN(n687) );
  XOR2_X1 U772 ( .A(n687), .B(KEYINPUT26), .Z(n689) );
  NAND2_X1 U773 ( .A1(n733), .A2(G1341), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U775 ( .A1(n1016), .A2(n690), .ZN(n692) );
  NOR2_X1 U776 ( .A1(n692), .A2(n1001), .ZN(n691) );
  XNOR2_X1 U777 ( .A(n691), .B(KEYINPUT103), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n692), .A2(n1001), .ZN(n696) );
  INV_X1 U779 ( .A(n720), .ZN(n699) );
  BUF_X1 U780 ( .A(n699), .Z(n715) );
  NOR2_X1 U781 ( .A1(n715), .A2(G1348), .ZN(n694) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n733), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n707) );
  INV_X1 U786 ( .A(KEYINPUT104), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n699), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  XOR2_X1 U789 ( .A(G1956), .B(KEYINPUT100), .Z(n918) );
  NOR2_X1 U790 ( .A1(n699), .A2(n918), .ZN(n701) );
  NOR2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT101), .ZN(n708) );
  XNOR2_X1 U793 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n707), .A2(n706), .ZN(n712) );
  NAND2_X1 U795 ( .A1(n708), .A2(G299), .ZN(n710) );
  XNOR2_X1 U796 ( .A(KEYINPUT102), .B(KEYINPUT28), .ZN(n709) );
  XNOR2_X1 U797 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U799 ( .A(n714), .B(n713), .ZN(n719) );
  INV_X1 U800 ( .A(G1961), .ZN(n930) );
  NAND2_X1 U801 ( .A1(n733), .A2(n930), .ZN(n717) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U803 ( .A1(n715), .A2(n945), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n725) );
  NAND2_X1 U805 ( .A1(n725), .A2(G171), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n732) );
  NAND2_X1 U807 ( .A1(G8), .A2(n720), .ZN(n778) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n778), .ZN(n747) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n733), .ZN(n744) );
  NOR2_X1 U810 ( .A1(n747), .A2(n744), .ZN(n721) );
  NAND2_X1 U811 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n722), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G168), .A2(n723), .ZN(n724) );
  XNOR2_X1 U814 ( .A(n724), .B(KEYINPUT105), .ZN(n727) );
  OR2_X1 U815 ( .A1(n725), .A2(G171), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n730) );
  XOR2_X1 U817 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n728) );
  XNOR2_X1 U818 ( .A(KEYINPUT31), .B(n728), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n745) );
  NAND2_X1 U821 ( .A1(n745), .A2(G286), .ZN(n739) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n778), .ZN(n735) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U825 ( .A1(n736), .A2(G303), .ZN(n737) );
  XNOR2_X1 U826 ( .A(n737), .B(KEYINPUT108), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U828 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U830 ( .A(KEYINPUT32), .B(n743), .ZN(n767) );
  NAND2_X1 U831 ( .A1(G8), .A2(n744), .ZN(n749) );
  INV_X1 U832 ( .A(n745), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n765) );
  NAND2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  INV_X1 U836 ( .A(n778), .ZN(n770) );
  NAND2_X1 U837 ( .A1(n1004), .A2(n770), .ZN(n757) );
  INV_X1 U838 ( .A(n757), .ZN(n750) );
  AND2_X1 U839 ( .A1(n765), .A2(n750), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n756), .A2(KEYINPUT33), .ZN(n751) );
  OR2_X1 U842 ( .A1(n751), .A2(n778), .ZN(n761) );
  AND2_X1 U843 ( .A1(n752), .A2(n761), .ZN(n753) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n1009) );
  AND2_X1 U845 ( .A1(n753), .A2(n1009), .ZN(n754) );
  AND2_X1 U846 ( .A1(n767), .A2(n754), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n1019) );
  OR2_X1 U849 ( .A1(n757), .A2(n1019), .ZN(n759) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n760) );
  AND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U853 ( .A1(n1009), .A2(n762), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n774) );
  AND2_X1 U855 ( .A1(n765), .A2(n778), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n772) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n768) );
  NAND2_X1 U858 ( .A1(G8), .A2(n768), .ZN(n769) );
  OR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT110), .ZN(n781) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U864 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U866 ( .A(KEYINPUT99), .B(n779), .Z(n780) );
  NOR2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n812) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n827) );
  XNOR2_X1 U869 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G128), .A2(n882), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G116), .A2(n883), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT35), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n788), .B(n787), .ZN(n793) );
  NAND2_X1 U875 ( .A1(G140), .A2(n886), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G104), .A2(n887), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n791), .ZN(n792) );
  NOR2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U880 ( .A(KEYINPUT36), .B(n794), .ZN(n872) );
  XNOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NOR2_X1 U882 ( .A1(n872), .A2(n825), .ZN(n991) );
  NAND2_X1 U883 ( .A1(n827), .A2(n991), .ZN(n822) );
  NAND2_X1 U884 ( .A1(G107), .A2(n883), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(KEYINPUT98), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G131), .A2(n886), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G95), .A2(n887), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G119), .A2(n882), .ZN(n798) );
  XNOR2_X1 U890 ( .A(KEYINPUT97), .B(n798), .ZN(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n876) );
  AND2_X1 U893 ( .A1(n876), .A2(G1991), .ZN(n975) );
  NAND2_X1 U894 ( .A1(G117), .A2(n883), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G141), .A2(n886), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n887), .A2(G105), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n882), .A2(G129), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n877) );
  AND2_X1 U902 ( .A1(n877), .A2(G1996), .ZN(n979) );
  OR2_X1 U903 ( .A1(n975), .A2(n979), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n810), .A2(n827), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n822), .A2(n816), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n814) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n1018) );
  NAND2_X1 U908 ( .A1(n1018), .A2(n827), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n830) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n877), .ZN(n815) );
  XOR2_X1 U911 ( .A(KEYINPUT111), .B(n815), .Z(n983) );
  INV_X1 U912 ( .A(n816), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n876), .ZN(n974) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n974), .A2(n817), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n983), .A2(n820), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n824), .B(KEYINPUT112), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n872), .A2(n825), .ZN(n988) );
  NAND2_X1 U922 ( .A1(n826), .A2(n988), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U925 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U928 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G188) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G325) );
  XNOR2_X1 U932 ( .A(KEYINPUT113), .B(G325), .ZN(G261) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  XOR2_X1 U937 ( .A(G2096), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2678), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n840), .B(KEYINPUT114), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2090), .B(G2072), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2100), .Z(n844) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1981), .Z(n848) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1971), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n849), .B(KEYINPUT41), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U953 ( .A(G2474), .B(G1956), .Z(n853) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1961), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G112), .A2(n883), .ZN(n857) );
  NAND2_X1 U958 ( .A1(G136), .A2(n886), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U960 ( .A1(G124), .A2(n882), .ZN(n858) );
  XOR2_X1 U961 ( .A(KEYINPUT115), .B(n858), .Z(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G100), .A2(n887), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G139), .A2(n886), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G103), .A2(n887), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G127), .A2(n882), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G115), .A2(n883), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n868), .Z(n869) );
  NOR2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n970) );
  XOR2_X1 U974 ( .A(G160), .B(n970), .Z(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n881) );
  XOR2_X1 U976 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n874) );
  XNOR2_X1 U977 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U978 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U979 ( .A(n875), .B(G162), .Z(n879) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U982 ( .A(n881), .B(n880), .Z(n895) );
  NAND2_X1 U983 ( .A1(G130), .A2(n882), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G118), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G142), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n981), .B(n893), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n896), .B(G164), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n1016), .B(G286), .ZN(n901) );
  XNOR2_X1 U996 ( .A(G301), .B(n1001), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n904) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n910) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n911) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n911), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(n917), .A2(G319), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n917), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(n918), .B(G20), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G19), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(G6), .B(G1981), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT59), .B(G1348), .Z(n923) );
  XNOR2_X1 U1025 ( .A(G4), .B(n923), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1027 ( .A(KEYINPUT60), .B(n926), .Z(n928) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G21), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT126), .B(n929), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n930), .B(G5), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n940) );
  XOR2_X1 U1033 ( .A(G1986), .B(G24), .Z(n936) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1038 ( .A(KEYINPUT58), .B(n937), .Z(n938) );
  XNOR2_X1 U1039 ( .A(KEYINPUT127), .B(n938), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n941), .Z(n942) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n942), .ZN(n969) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n996) );
  XOR2_X1 U1044 ( .A(KEYINPUT124), .B(G34), .Z(n944) );
  XNOR2_X1 U1045 ( .A(G2084), .B(KEYINPUT54), .ZN(n943) );
  XNOR2_X1 U1046 ( .A(n944), .B(n943), .ZN(n963) );
  XNOR2_X1 U1047 ( .A(G2090), .B(G35), .ZN(n961) );
  XNOR2_X1 U1048 ( .A(G27), .B(n945), .ZN(n949) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1051 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1053 ( .A(G32), .B(G1996), .Z(n950) );
  XNOR2_X1 U1054 ( .A(KEYINPUT121), .B(n950), .ZN(n951) );
  NOR2_X1 U1055 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1056 ( .A(KEYINPUT122), .B(n953), .ZN(n957) );
  XOR2_X1 U1057 ( .A(G25), .B(G1991), .Z(n954) );
  NAND2_X1 U1058 ( .A1(n954), .A2(G28), .ZN(n955) );
  XOR2_X1 U1059 ( .A(KEYINPUT120), .B(n955), .Z(n956) );
  NAND2_X1 U1060 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1061 ( .A(n958), .B(KEYINPUT123), .ZN(n959) );
  XNOR2_X1 U1062 ( .A(n959), .B(KEYINPUT53), .ZN(n960) );
  NOR2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1065 ( .A(n996), .B(n964), .ZN(n966) );
  INV_X1 U1066 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1067 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n967), .ZN(n968) );
  NOR2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n1000) );
  XOR2_X1 U1070 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1071 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1073 ( .A(KEYINPUT50), .B(n973), .Z(n994) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1081 ( .A(KEYINPUT118), .B(n984), .Z(n985) );
  XOR2_X1 U1082 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT119), .B(n992), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT52), .B(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(G29), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  XOR2_X1 U1092 ( .A(G16), .B(KEYINPUT56), .Z(n1024) );
  XNOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT125), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(n1001), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(G1971), .A2(G303), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(G1956), .B(G299), .Z(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G168), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1103 ( .A(KEYINPUT57), .B(n1011), .Z(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G1341), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1027), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

