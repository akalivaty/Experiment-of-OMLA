

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731;

  NAND2_X1 U367 ( .A1(n346), .A2(n601), .ZN(n402) );
  NOR2_X1 U368 ( .A1(n687), .A2(n345), .ZN(n346) );
  INV_X1 U369 ( .A(KEYINPUT79), .ZN(n345) );
  INV_X1 U370 ( .A(n686), .ZN(n356) );
  AND2_X1 U371 ( .A1(n608), .A2(n576), .ZN(n577) );
  XNOR2_X1 U372 ( .A(n572), .B(n571), .ZN(n608) );
  AND2_X1 U373 ( .A1(n506), .A2(n378), .ZN(n650) );
  AND2_X1 U374 ( .A1(n562), .A2(n587), .ZN(n569) );
  NOR2_X1 U375 ( .A1(n670), .A2(n669), .ZN(n533) );
  BUF_X1 U376 ( .A(n380), .Z(n378) );
  NOR2_X1 U377 ( .A1(n653), .A2(n563), .ZN(n656) );
  NOR2_X1 U378 ( .A1(G902), .A2(n693), .ZN(n504) );
  XNOR2_X1 U379 ( .A(n468), .B(n467), .ZN(n653) );
  XNOR2_X1 U380 ( .A(n418), .B(KEYINPUT68), .ZN(n718) );
  XNOR2_X1 U381 ( .A(n417), .B(G146), .ZN(n484) );
  XNOR2_X1 U382 ( .A(n440), .B(n441), .ZN(n443) );
  INV_X1 U383 ( .A(G953), .ZN(n706) );
  OR2_X2 U384 ( .A1(n505), .A2(n379), .ZN(n561) );
  NOR2_X2 U385 ( .A1(n579), .A2(n587), .ZN(n371) );
  XNOR2_X2 U386 ( .A(n400), .B(KEYINPUT74), .ZN(n579) );
  XNOR2_X2 U387 ( .A(n504), .B(n401), .ZN(n522) );
  INV_X1 U388 ( .A(G469), .ZN(n401) );
  NOR2_X1 U389 ( .A1(n534), .A2(n554), .ZN(n516) );
  XNOR2_X1 U390 ( .A(n556), .B(n555), .ZN(n583) );
  XNOR2_X1 U391 ( .A(n444), .B(G472), .ZN(n573) );
  XNOR2_X1 U392 ( .A(n443), .B(n442), .ZN(n496) );
  XNOR2_X1 U393 ( .A(n422), .B(G143), .ZN(n483) );
  XNOR2_X1 U394 ( .A(n485), .B(G137), .ZN(n440) );
  INV_X1 U395 ( .A(G128), .ZN(n422) );
  INV_X1 U396 ( .A(G125), .ZN(n417) );
  XOR2_X1 U397 ( .A(G134), .B(n483), .Z(n442) );
  NAND2_X1 U398 ( .A1(n546), .A2(n545), .ZN(n603) );
  XNOR2_X1 U399 ( .A(n384), .B(n383), .ZN(n546) );
  INV_X1 U400 ( .A(KEYINPUT48), .ZN(n383) );
  NOR2_X1 U401 ( .A1(n587), .A2(n474), .ZN(n395) );
  XNOR2_X1 U402 ( .A(n434), .B(n433), .ZN(n479) );
  XNOR2_X1 U403 ( .A(G101), .B(KEYINPUT3), .ZN(n433) );
  INV_X1 U404 ( .A(G119), .ZN(n431) );
  INV_X1 U405 ( .A(KEYINPUT84), .ZN(n391) );
  NAND2_X1 U406 ( .A1(n388), .A2(n387), .ZN(n386) );
  XOR2_X1 U407 ( .A(KEYINPUT78), .B(KEYINPUT8), .Z(n428) );
  XNOR2_X1 U408 ( .A(n482), .B(KEYINPUT87), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n522), .B(KEYINPUT1), .ZN(n380) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n435) );
  XNOR2_X1 U411 ( .A(n437), .B(G146), .ZN(n438) );
  XOR2_X1 U412 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n437) );
  INV_X1 U413 ( .A(n439), .ZN(n441) );
  XNOR2_X1 U414 ( .A(KEYINPUT16), .B(G122), .ZN(n478) );
  XNOR2_X1 U415 ( .A(n355), .B(n456), .ZN(n457) );
  XNOR2_X1 U416 ( .A(n495), .B(n455), .ZN(n355) );
  INV_X1 U417 ( .A(n442), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n425) );
  XNOR2_X1 U419 ( .A(KEYINPUT100), .B(KEYINPUT7), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n423), .B(KEYINPUT101), .ZN(n364) );
  XNOR2_X1 U421 ( .A(G122), .B(KEYINPUT9), .ZN(n423) );
  NAND2_X1 U422 ( .A1(n382), .A2(KEYINPUT2), .ZN(n381) );
  INV_X1 U423 ( .A(n603), .ZN(n382) );
  NOR2_X1 U424 ( .A1(n640), .A2(n513), .ZN(n392) );
  XNOR2_X1 U425 ( .A(n370), .B(n399), .ZN(n398) );
  INV_X1 U426 ( .A(KEYINPUT34), .ZN(n399) );
  XNOR2_X1 U427 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U428 ( .A(n430), .B(G478), .ZN(n531) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n430) );
  INV_X1 U430 ( .A(KEYINPUT102), .ZN(n359) );
  OR2_X1 U431 ( .A1(n698), .A2(G902), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n568), .B(n567), .ZN(n590) );
  NAND2_X1 U433 ( .A1(n692), .A2(G475), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT86), .B(n607), .Z(n691) );
  NOR2_X1 U435 ( .A1(n378), .A2(n656), .ZN(n657) );
  XNOR2_X1 U436 ( .A(n386), .B(n540), .ZN(n385) );
  XOR2_X1 U437 ( .A(KEYINPUT21), .B(n473), .Z(n654) );
  XNOR2_X1 U438 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U439 ( .A(G116), .B(G113), .ZN(n432) );
  XOR2_X1 U440 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n455) );
  XNOR2_X1 U441 ( .A(G143), .B(G122), .ZN(n411) );
  XOR2_X1 U442 ( .A(KEYINPUT12), .B(G140), .Z(n412) );
  INV_X1 U443 ( .A(KEYINPUT2), .ZN(n406) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n446) );
  INV_X1 U445 ( .A(G237), .ZN(n475) );
  AND2_X1 U446 ( .A1(n469), .A2(n653), .ZN(n508) );
  INV_X1 U447 ( .A(KEYINPUT109), .ZN(n509) );
  INV_X1 U448 ( .A(G902), .ZN(n476) );
  XNOR2_X1 U449 ( .A(n496), .B(n495), .ZN(n719) );
  XOR2_X1 U450 ( .A(G101), .B(G146), .Z(n498) );
  XNOR2_X1 U451 ( .A(G110), .B(G107), .ZN(n477) );
  XNOR2_X1 U452 ( .A(n481), .B(n353), .ZN(n488) );
  OR2_X1 U453 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U454 ( .A(n496), .B(n396), .ZN(n611) );
  XNOR2_X1 U455 ( .A(n479), .B(n397), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n438), .B(n436), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n457), .B(n718), .ZN(n462) );
  XNOR2_X1 U458 ( .A(G119), .B(G137), .ZN(n459) );
  XNOR2_X1 U459 ( .A(n426), .B(n361), .ZN(n698) );
  XNOR2_X1 U460 ( .A(n429), .B(n362), .ZN(n361) );
  XNOR2_X1 U461 ( .A(G116), .B(G107), .ZN(n424) );
  XNOR2_X1 U462 ( .A(n689), .B(n369), .ZN(n368) );
  INV_X1 U463 ( .A(KEYINPUT80), .ZN(n369) );
  NOR2_X1 U464 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U465 ( .A1(n542), .A2(n378), .ZN(n543) );
  XNOR2_X1 U466 ( .A(n560), .B(n559), .ZN(n728) );
  NAND2_X1 U467 ( .A1(n398), .A2(n557), .ZN(n560) );
  AND2_X1 U468 ( .A1(n505), .A2(n379), .ZN(n588) );
  INV_X1 U469 ( .A(KEYINPUT60), .ZN(n372) );
  NAND2_X1 U470 ( .A1(n374), .A2(n691), .ZN(n373) );
  XNOR2_X1 U471 ( .A(n375), .B(n606), .ZN(n374) );
  XNOR2_X1 U472 ( .A(n366), .B(n365), .ZN(G75) );
  INV_X1 U473 ( .A(KEYINPUT53), .ZN(n365) );
  NAND2_X1 U474 ( .A1(n368), .A2(n367), .ZN(n366) );
  AND2_X1 U475 ( .A1(n690), .A2(n706), .ZN(n367) );
  XOR2_X1 U476 ( .A(n544), .B(n529), .Z(n347) );
  XNOR2_X1 U477 ( .A(G140), .B(KEYINPUT70), .ZN(n495) );
  XNOR2_X1 U478 ( .A(n493), .B(n492), .ZN(n544) );
  INV_X1 U479 ( .A(n544), .ZN(n354) );
  AND2_X1 U480 ( .A1(n357), .A2(n356), .ZN(n348) );
  XOR2_X1 U481 ( .A(n543), .B(KEYINPUT43), .Z(n349) );
  AND2_X1 U482 ( .A1(n528), .A2(n527), .ZN(n350) );
  XNOR2_X1 U483 ( .A(n719), .B(n503), .ZN(n693) );
  AND2_X1 U484 ( .A1(n578), .A2(KEYINPUT72), .ZN(n351) );
  XNOR2_X1 U485 ( .A(n352), .B(n351), .ZN(n595) );
  NAND2_X1 U486 ( .A1(n577), .A2(n728), .ZN(n352) );
  NAND2_X1 U487 ( .A1(n354), .A2(n667), .ZN(n515) );
  NAND2_X1 U488 ( .A1(n404), .A2(n376), .ZN(n403) );
  NAND2_X1 U489 ( .A1(n598), .A2(n356), .ZN(n377) );
  NOR2_X1 U490 ( .A1(n358), .A2(n599), .ZN(n600) );
  INV_X1 U491 ( .A(n358), .ZN(n357) );
  NOR2_X1 U492 ( .A1(n358), .A2(KEYINPUT79), .ZN(n598) );
  XNOR2_X1 U493 ( .A(n358), .B(n720), .ZN(n721) );
  XNOR2_X2 U494 ( .A(n603), .B(n547), .ZN(n358) );
  NAND2_X1 U495 ( .A1(n674), .A2(n583), .ZN(n370) );
  XNOR2_X1 U496 ( .A(n371), .B(n548), .ZN(n674) );
  XNOR2_X1 U497 ( .A(n373), .B(n372), .ZN(G60) );
  NAND2_X1 U498 ( .A1(n377), .A2(n406), .ZN(n376) );
  NAND2_X1 U499 ( .A1(n656), .A2(n380), .ZN(n400) );
  INV_X1 U500 ( .A(n378), .ZN(n505) );
  INV_X1 U501 ( .A(n653), .ZN(n379) );
  XNOR2_X2 U502 ( .A(n538), .B(KEYINPUT39), .ZN(n541) );
  AND2_X2 U503 ( .A1(n541), .A2(n643), .ZN(n539) );
  XNOR2_X2 U504 ( .A(n539), .B(KEYINPUT40), .ZN(n730) );
  XNOR2_X2 U505 ( .A(n597), .B(n596), .ZN(n686) );
  XNOR2_X2 U506 ( .A(G902), .B(KEYINPUT15), .ZN(n599) );
  NOR2_X2 U507 ( .A1(n686), .A2(n381), .ZN(n687) );
  NAND2_X1 U508 ( .A1(n389), .A2(n385), .ZN(n384) );
  INV_X1 U509 ( .A(n731), .ZN(n387) );
  INV_X1 U510 ( .A(n730), .ZN(n388) );
  AND2_X1 U511 ( .A1(n390), .A2(n350), .ZN(n389) );
  XNOR2_X1 U512 ( .A(n650), .B(n391), .ZN(n390) );
  NAND2_X1 U513 ( .A1(n393), .A2(n392), .ZN(n542) );
  XNOR2_X1 U514 ( .A(n395), .B(n394), .ZN(n393) );
  INV_X1 U515 ( .A(KEYINPUT107), .ZN(n394) );
  NAND2_X2 U516 ( .A1(n402), .A2(n403), .ZN(n692) );
  NOR2_X1 U517 ( .A1(n687), .A2(n599), .ZN(n404) );
  XNOR2_X1 U518 ( .A(n696), .B(n695), .ZN(n697) );
  AND2_X1 U519 ( .A1(n594), .A2(n593), .ZN(n407) );
  INV_X1 U520 ( .A(n638), .ZN(n527) );
  INV_X1 U521 ( .A(KEYINPUT46), .ZN(n540) );
  XNOR2_X1 U522 ( .A(n509), .B(KEYINPUT28), .ZN(n510) );
  XNOR2_X1 U523 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n693), .B(n694), .ZN(n695) );
  XNOR2_X1 U525 ( .A(KEYINPUT13), .B(G475), .ZN(n421) );
  XOR2_X1 U526 ( .A(KEYINPUT69), .B(G131), .Z(n439) );
  XNOR2_X1 U527 ( .A(n439), .B(G113), .ZN(n408) );
  XNOR2_X1 U528 ( .A(n408), .B(G104), .ZN(n416) );
  XOR2_X1 U529 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n410) );
  NAND2_X1 U530 ( .A1(G214), .A2(n435), .ZN(n409) );
  XNOR2_X1 U531 ( .A(n410), .B(n409), .ZN(n414) );
  XNOR2_X1 U532 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U533 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U534 ( .A(n416), .B(n415), .Z(n419) );
  XNOR2_X1 U535 ( .A(n484), .B(KEYINPUT10), .ZN(n418) );
  XNOR2_X1 U536 ( .A(n419), .B(n718), .ZN(n605) );
  NOR2_X1 U537 ( .A1(G902), .A2(n605), .ZN(n420) );
  XNOR2_X1 U538 ( .A(n421), .B(n420), .ZN(n525) );
  XNOR2_X1 U539 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U540 ( .A1(G234), .A2(n706), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n428), .B(n427), .ZN(n458) );
  NAND2_X1 U542 ( .A1(G217), .A2(n458), .ZN(n429) );
  NAND2_X1 U543 ( .A1(n525), .A2(n531), .ZN(n640) );
  XNOR2_X1 U544 ( .A(n432), .B(n431), .ZN(n434) );
  AND2_X1 U545 ( .A1(n435), .A2(G210), .ZN(n436) );
  XOR2_X2 U546 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n485) );
  NAND2_X1 U547 ( .A1(n611), .A2(n476), .ZN(n444) );
  INV_X1 U548 ( .A(n573), .ZN(n581) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n445) );
  XNOR2_X1 U550 ( .A(n581), .B(n445), .ZN(n587) );
  XNOR2_X1 U551 ( .A(n446), .B(KEYINPUT14), .ZN(n448) );
  NAND2_X1 U552 ( .A1(n448), .A2(G952), .ZN(n447) );
  XOR2_X1 U553 ( .A(KEYINPUT89), .B(n447), .Z(n681) );
  NOR2_X1 U554 ( .A1(G953), .A2(n681), .ZN(n551) );
  NAND2_X1 U555 ( .A1(n448), .A2(G902), .ZN(n449) );
  XOR2_X1 U556 ( .A(KEYINPUT90), .B(n449), .Z(n549) );
  NAND2_X1 U557 ( .A1(G953), .A2(n549), .ZN(n450) );
  NOR2_X1 U558 ( .A1(G900), .A2(n450), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n451), .B(KEYINPUT106), .ZN(n452) );
  NOR2_X1 U560 ( .A1(n551), .A2(n452), .ZN(n521) );
  INV_X1 U561 ( .A(n521), .ZN(n469) );
  XOR2_X1 U562 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n454) );
  XNOR2_X1 U563 ( .A(G128), .B(G110), .ZN(n453) );
  XNOR2_X1 U564 ( .A(n454), .B(n453), .ZN(n456) );
  NAND2_X1 U565 ( .A1(G221), .A2(n458), .ZN(n460) );
  XNOR2_X1 U566 ( .A(n462), .B(n461), .ZN(n703) );
  NOR2_X1 U567 ( .A1(G902), .A2(n703), .ZN(n468) );
  NAND2_X1 U568 ( .A1(n599), .A2(G234), .ZN(n463) );
  XNOR2_X1 U569 ( .A(n463), .B(KEYINPUT94), .ZN(n464) );
  XNOR2_X1 U570 ( .A(KEYINPUT20), .B(n464), .ZN(n470) );
  NAND2_X1 U571 ( .A1(G217), .A2(n470), .ZN(n466) );
  INV_X1 U572 ( .A(KEYINPUT25), .ZN(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n472) );
  NAND2_X1 U574 ( .A1(G221), .A2(n470), .ZN(n471) );
  NAND2_X1 U575 ( .A1(n508), .A2(n654), .ZN(n474) );
  NAND2_X1 U576 ( .A1(n476), .A2(n475), .ZN(n490) );
  NAND2_X1 U577 ( .A1(n490), .A2(G214), .ZN(n667) );
  XNOR2_X1 U578 ( .A(n477), .B(G104), .ZN(n500) );
  XNOR2_X1 U579 ( .A(n500), .B(n478), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n480), .B(n479), .ZN(n712) );
  NAND2_X1 U581 ( .A1(n706), .A2(G224), .ZN(n481) );
  XNOR2_X1 U582 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n486) );
  XNOR2_X1 U584 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n712), .B(n489), .ZN(n617) );
  NAND2_X1 U587 ( .A1(n617), .A2(n599), .ZN(n493) );
  NAND2_X1 U588 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U589 ( .A(n491), .B(KEYINPUT88), .ZN(n492) );
  NOR2_X1 U590 ( .A1(n542), .A2(n544), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n494), .B(KEYINPUT36), .ZN(n506) );
  NAND2_X1 U592 ( .A1(G227), .A2(n706), .ZN(n497) );
  XNOR2_X1 U593 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U594 ( .A(n499), .B(KEYINPUT75), .Z(n502) );
  XNOR2_X1 U595 ( .A(n500), .B(KEYINPUT76), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U597 ( .A1(n525), .A2(n531), .ZN(n646) );
  INV_X1 U598 ( .A(n640), .ZN(n643) );
  OR2_X1 U599 ( .A1(n646), .A2(n643), .ZN(n585) );
  INV_X1 U600 ( .A(n585), .ZN(n671) );
  INV_X1 U601 ( .A(n654), .ZN(n563) );
  NOR2_X1 U602 ( .A1(n563), .A2(n581), .ZN(n507) );
  AND2_X1 U603 ( .A1(n508), .A2(n507), .ZN(n511) );
  XNOR2_X1 U604 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U605 ( .A1(n512), .A2(n522), .ZN(n534) );
  INV_X1 U606 ( .A(n667), .ZN(n513) );
  XNOR2_X1 U607 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n514) );
  XNOR2_X1 U608 ( .A(n515), .B(n514), .ZN(n554) );
  XNOR2_X1 U609 ( .A(n516), .B(KEYINPUT77), .ZN(n639) );
  NOR2_X1 U610 ( .A1(n671), .A2(n639), .ZN(n517) );
  XNOR2_X1 U611 ( .A(n517), .B(KEYINPUT47), .ZN(n528) );
  XOR2_X1 U612 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n519) );
  NAND2_X1 U613 ( .A1(n573), .A2(n667), .ZN(n518) );
  XOR2_X1 U614 ( .A(n519), .B(n518), .Z(n520) );
  NOR2_X1 U615 ( .A1(n521), .A2(n520), .ZN(n524) );
  NAND2_X1 U616 ( .A1(n656), .A2(n522), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n523), .B(KEYINPUT97), .ZN(n582) );
  NAND2_X1 U618 ( .A1(n524), .A2(n582), .ZN(n536) );
  INV_X1 U619 ( .A(n525), .ZN(n530) );
  NOR2_X1 U620 ( .A1(n531), .A2(n530), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n557), .A2(n354), .ZN(n526) );
  NOR2_X1 U622 ( .A1(n536), .A2(n526), .ZN(n638) );
  XNOR2_X1 U623 ( .A(KEYINPUT73), .B(KEYINPUT38), .ZN(n529) );
  NAND2_X1 U624 ( .A1(n347), .A2(n667), .ZN(n670) );
  NAND2_X1 U625 ( .A1(n531), .A2(n530), .ZN(n669) );
  XNOR2_X1 U626 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n533), .B(n532), .ZN(n683) );
  NOR2_X1 U628 ( .A1(n534), .A2(n683), .ZN(n535) );
  XNOR2_X1 U629 ( .A(n535), .B(KEYINPUT42), .ZN(n731) );
  INV_X1 U630 ( .A(n536), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n537), .A2(n347), .ZN(n538) );
  NAND2_X1 U632 ( .A1(n541), .A2(n646), .ZN(n652) );
  NAND2_X1 U633 ( .A1(n349), .A2(n544), .ZN(n609) );
  AND2_X1 U634 ( .A1(n652), .A2(n609), .ZN(n545) );
  INV_X1 U635 ( .A(KEYINPUT81), .ZN(n547) );
  XNOR2_X1 U636 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n548) );
  NOR2_X1 U637 ( .A1(G898), .A2(n706), .ZN(n713) );
  AND2_X1 U638 ( .A1(n713), .A2(n549), .ZN(n550) );
  OR2_X1 U639 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U640 ( .A(n552), .B(KEYINPUT91), .ZN(n553) );
  INV_X1 U641 ( .A(KEYINPUT0), .ZN(n555) );
  INV_X1 U642 ( .A(KEYINPUT82), .ZN(n558) );
  XNOR2_X1 U643 ( .A(n558), .B(KEYINPUT35), .ZN(n559) );
  XNOR2_X1 U644 ( .A(n561), .B(KEYINPUT105), .ZN(n562) );
  NOR2_X1 U645 ( .A1(n669), .A2(n563), .ZN(n564) );
  XNOR2_X1 U646 ( .A(n564), .B(KEYINPUT104), .ZN(n565) );
  NAND2_X1 U647 ( .A1(n565), .A2(n583), .ZN(n568) );
  INV_X1 U648 ( .A(KEYINPUT66), .ZN(n566) );
  XNOR2_X1 U649 ( .A(n566), .B(KEYINPUT22), .ZN(n567) );
  NAND2_X1 U650 ( .A1(n569), .A2(n590), .ZN(n572) );
  INV_X1 U651 ( .A(KEYINPUT65), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n570), .B(KEYINPUT32), .ZN(n571) );
  NOR2_X1 U653 ( .A1(n378), .A2(n573), .ZN(n574) );
  AND2_X1 U654 ( .A1(n653), .A2(n574), .ZN(n575) );
  AND2_X1 U655 ( .A1(n590), .A2(n575), .ZN(n633) );
  INV_X1 U656 ( .A(n633), .ZN(n576) );
  INV_X1 U657 ( .A(KEYINPUT44), .ZN(n578) );
  NOR2_X1 U658 ( .A1(n579), .A2(n581), .ZN(n663) );
  NAND2_X1 U659 ( .A1(n663), .A2(n583), .ZN(n580) );
  XNOR2_X1 U660 ( .A(n580), .B(KEYINPUT31), .ZN(n647) );
  AND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n584) );
  AND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n630) );
  OR2_X1 U663 ( .A1(n647), .A2(n630), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n594) );
  AND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U666 ( .A1(n590), .A2(n589), .ZN(n623) );
  INV_X1 U667 ( .A(KEYINPUT72), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n591), .A2(KEYINPUT44), .ZN(n592) );
  AND2_X1 U669 ( .A1(n623), .A2(n592), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n595), .A2(n407), .ZN(n597) );
  INV_X1 U671 ( .A(KEYINPUT45), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n600), .A2(n356), .ZN(n601) );
  XOR2_X1 U673 ( .A(KEYINPUT85), .B(KEYINPUT59), .Z(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n706), .A2(G952), .ZN(n607) );
  XNOR2_X1 U676 ( .A(n608), .B(G119), .ZN(G21) );
  XNOR2_X1 U677 ( .A(n609), .B(G140), .ZN(G42) );
  NAND2_X1 U678 ( .A1(n692), .A2(G472), .ZN(n613) );
  XOR2_X1 U679 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n610) );
  XNOR2_X1 U680 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U682 ( .A1(n614), .A2(n691), .ZN(n615) );
  XNOR2_X1 U683 ( .A(n615), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U684 ( .A1(n692), .A2(G210), .ZN(n619) );
  XOR2_X1 U685 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n616) );
  XNOR2_X1 U686 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U687 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n620), .A2(n691), .ZN(n622) );
  XNOR2_X1 U689 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n622), .B(n621), .ZN(G51) );
  XNOR2_X1 U691 ( .A(G101), .B(KEYINPUT112), .ZN(n624) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(G3) );
  XOR2_X1 U693 ( .A(G104), .B(KEYINPUT113), .Z(n626) );
  NAND2_X1 U694 ( .A1(n630), .A2(n643), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n628) );
  XNOR2_X1 U697 ( .A(G107), .B(KEYINPUT114), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n629) );
  XOR2_X1 U699 ( .A(KEYINPUT26), .B(n629), .Z(n632) );
  NAND2_X1 U700 ( .A1(n630), .A2(n646), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(G9) );
  XOR2_X1 U702 ( .A(G110), .B(n633), .Z(G12) );
  INV_X1 U703 ( .A(n646), .ZN(n634) );
  NOR2_X1 U704 ( .A1(n634), .A2(n639), .ZN(n636) );
  XNOR2_X1 U705 ( .A(KEYINPUT29), .B(KEYINPUT116), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(G128), .B(n637), .ZN(G30) );
  XOR2_X1 U708 ( .A(G143), .B(n638), .Z(G45) );
  NOR2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U710 ( .A(G146), .B(KEYINPUT117), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(G48) );
  NAND2_X1 U712 ( .A1(n647), .A2(n643), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT118), .ZN(n645) );
  XNOR2_X1 U714 ( .A(G113), .B(n645), .ZN(G15) );
  XOR2_X1 U715 ( .A(G116), .B(KEYINPUT119), .Z(n649) );
  NAND2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(n648), .ZN(G18) );
  XNOR2_X1 U718 ( .A(G125), .B(n650), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n651), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U720 ( .A(G134), .B(n652), .ZN(G36) );
  NOR2_X1 U721 ( .A1(n654), .A2(n379), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT49), .B(n655), .ZN(n660) );
  XOR2_X1 U723 ( .A(KEYINPUT50), .B(n657), .Z(n658) );
  XNOR2_X1 U724 ( .A(KEYINPUT120), .B(n658), .ZN(n659) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n573), .A2(n661), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(KEYINPUT121), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT51), .B(n665), .ZN(n666) );
  NOR2_X1 U730 ( .A1(n683), .A2(n666), .ZN(n678) );
  NOR2_X1 U731 ( .A1(n347), .A2(n667), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n675) );
  INV_X1 U735 ( .A(n674), .ZN(n682) );
  NOR2_X1 U736 ( .A1(n675), .A2(n682), .ZN(n676) );
  XNOR2_X1 U737 ( .A(n676), .B(KEYINPUT122), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U739 ( .A(n679), .B(KEYINPUT52), .ZN(n680) );
  NOR2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U743 ( .A1(n348), .A2(KEYINPUT2), .ZN(n688) );
  INV_X1 U744 ( .A(n691), .ZN(n705) );
  BUF_X2 U745 ( .A(n692), .Z(n701) );
  NAND2_X1 U746 ( .A1(n701), .A2(G469), .ZN(n696) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  NOR2_X1 U748 ( .A1(n705), .A2(n697), .ZN(G54) );
  NAND2_X1 U749 ( .A1(n701), .A2(G478), .ZN(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n705), .A2(n700), .ZN(G63) );
  NAND2_X1 U752 ( .A1(n701), .A2(G217), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U754 ( .A1(n705), .A2(n704), .ZN(G66) );
  NAND2_X1 U755 ( .A1(n356), .A2(n706), .ZN(n711) );
  XOR2_X1 U756 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n708) );
  NAND2_X1 U757 ( .A1(G224), .A2(G953), .ZN(n707) );
  XNOR2_X1 U758 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U759 ( .A1(n709), .A2(G898), .ZN(n710) );
  NAND2_X1 U760 ( .A1(n711), .A2(n710), .ZN(n716) );
  INV_X1 U761 ( .A(n712), .ZN(n714) );
  NOR2_X1 U762 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U763 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U764 ( .A(KEYINPUT124), .B(n717), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n719), .B(n718), .ZN(n723) );
  INV_X1 U766 ( .A(n723), .ZN(n720) );
  NOR2_X1 U767 ( .A1(G953), .A2(n721), .ZN(n722) );
  XNOR2_X1 U768 ( .A(KEYINPUT125), .B(n722), .ZN(n727) );
  XNOR2_X1 U769 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U770 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n727), .A2(n726), .ZN(G72) );
  XNOR2_X1 U773 ( .A(n728), .B(G122), .ZN(n729) );
  XNOR2_X1 U774 ( .A(n729), .B(KEYINPUT126), .ZN(G24) );
  XOR2_X1 U775 ( .A(G131), .B(n730), .Z(G33) );
  XOR2_X1 U776 ( .A(G137), .B(n731), .Z(G39) );
endmodule

