//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G116), .A2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n201), .A2(new_n212), .B1(new_n202), .B2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n211), .B(new_n214), .C1(G107), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT66), .B(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT67), .B(G238), .Z(new_n218));
  OAI21_X1  g0018(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT68), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n207), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n226));
  AND3_X1   g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n207), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n223), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n213), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT70), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G223), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(G1698), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n260), .A2(G222), .B1(G77), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(KEYINPUT69), .B(G226), .Z(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n264), .A3(G274), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(G190), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n204), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n230), .A2(G33), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT71), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n229), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n283), .A2(new_n288), .B1(new_n201), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n288), .B1(new_n289), .B2(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT73), .B(G200), .Z(new_n297));
  AOI21_X1  g0097(.A(new_n264), .B1(new_n259), .B2(new_n261), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n274), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n276), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n276), .A2(new_n299), .A3(new_n296), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n281), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n279), .B1(G20), .B2(G77), .ZN(new_n306));
  INV_X1    g0106(.A(G87), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT15), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT72), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n306), .B1(new_n315), .B2(new_n282), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n288), .B1(new_n209), .B2(new_n291), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n293), .A2(G77), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n218), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n258), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n260), .A2(G232), .B1(G107), .B2(new_n255), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n264), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n270), .A2(G244), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n273), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n319), .B1(new_n326), .B2(new_n297), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n323), .A2(new_n325), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n330), .B1(new_n318), .B2(new_n317), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n323), .B2(new_n325), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n327), .A2(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n266), .A2(new_n330), .A3(new_n275), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(new_n298), .B2(new_n274), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n295), .A3(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n304), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n305), .A2(new_n290), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n293), .B2(new_n305), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n230), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n230), .A4(new_n344), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(KEYINPUT77), .A3(new_n346), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n216), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n280), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT66), .A2(G68), .ZN(new_n355));
  NOR2_X1   g0155(.A1(KEYINPUT66), .A2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(G58), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n224), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n354), .B1(new_n359), .B2(G20), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT16), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n255), .B2(new_n230), .ZN(new_n362));
  INV_X1    g0162(.A(new_n349), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n360), .A3(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n288), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n340), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n289), .B1(G41), .B2(G45), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n264), .A2(G232), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n368), .B1(new_n273), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(G223), .A2(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n212), .A2(G1698), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(new_n253), .C2(new_n254), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n264), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n273), .A2(new_n370), .A3(new_n368), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n372), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n273), .A2(new_n370), .A3(new_n368), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n382), .A2(new_n371), .A3(new_n377), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n383), .B2(G200), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT17), .B1(new_n367), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n352), .A2(new_n360), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n288), .ZN(new_n390));
  INV_X1    g0190(.A(new_n354), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n224), .B1(new_n216), .B2(G58), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n230), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n203), .B1(new_n347), .B2(new_n349), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n390), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n340), .A4(new_n384), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n386), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n340), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n389), .B2(new_n396), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n383), .A2(new_n332), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n382), .A2(new_n371), .A3(new_n377), .A4(new_n330), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT18), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n383), .A2(G179), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n332), .B2(new_n383), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n367), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n400), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n217), .A2(KEYINPUT12), .A3(new_n291), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n216), .A2(new_n230), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n280), .A2(new_n201), .B1(new_n282), .B2(new_n209), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n288), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n413), .B1(KEYINPUT12), .B2(new_n291), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n293), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n203), .B1(new_n419), .B2(KEYINPUT12), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n416), .A2(new_n417), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n273), .B(KEYINPUT74), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n270), .A2(G238), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n213), .A2(G1698), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G226), .B2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n255), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n265), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n426), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT13), .B1(new_n433), .B2(new_n423), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n422), .B1(new_n435), .B2(new_n379), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  INV_X1    g0237(.A(G200), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT75), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT75), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n440), .A3(G200), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n436), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n332), .B1(new_n432), .B2(new_n434), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n443), .A2(new_n444), .B1(new_n435), .B2(new_n330), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT76), .B1(new_n443), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n422), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n338), .A2(new_n412), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n338), .A2(KEYINPUT79), .A3(new_n412), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n350), .A2(G107), .A3(new_n351), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT6), .A3(G97), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n459), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n460), .B1(new_n464), .B2(KEYINPUT6), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n390), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n291), .A2(new_n461), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n284), .A2(new_n285), .B1(G1), .B2(G13), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n289), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n287), .A3(new_n290), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n461), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(G244), .C1(new_n254), .C2(new_n253), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n210), .B1(new_n343), .B2(new_n344), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n256), .B1(new_n479), .B2(KEYINPUT4), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n265), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n289), .B(G45), .C1(new_n267), .C2(KEYINPUT5), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n265), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n264), .A2(G274), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n485), .A2(G257), .B1(new_n486), .B2(new_n484), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n467), .A2(new_n472), .B1(new_n488), .B2(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT80), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n481), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(new_n332), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n467), .A2(new_n472), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(G200), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(G190), .A3(new_n492), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(KEYINPUT81), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n490), .A2(new_n500), .A3(G190), .A4(new_n492), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n494), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT84), .B1(new_n315), .B2(new_n471), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n290), .A2(new_n470), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n288), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT72), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT72), .B1(new_n308), .B2(new_n310), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n315), .A2(new_n291), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n230), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n230), .A2(G33), .A3(G97), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT82), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT19), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n230), .B1(new_n521), .B2(new_n427), .ZN(new_n522));
  OR2_X1    g0322(.A1(KEYINPUT83), .A2(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT83), .A2(G87), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n463), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n520), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n512), .B1(new_n526), .B2(new_n390), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT85), .B1(new_n511), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n520), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n427), .B1(new_n516), .B2(new_n518), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n525), .B1(new_n530), .B2(G20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n288), .B1(new_n291), .B2(new_n315), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n503), .A2(new_n510), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT85), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OR3_X1    g0336(.A1(new_n268), .A2(G1), .A3(G274), .ZN(new_n537));
  INV_X1    g0337(.A(G250), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n268), .B2(G1), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n264), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G116), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n342), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G238), .A2(G1698), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n210), .B2(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n343), .A2(new_n344), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(new_n264), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G169), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n330), .B2(new_n547), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n528), .A2(new_n536), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n390), .B1(new_n529), .B2(new_n531), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n508), .A2(new_n290), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n471), .A2(new_n307), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OR2_X1    g0354(.A1(G238), .A2(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n210), .A2(G1698), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n253), .C2(new_n254), .ZN(new_n557));
  INV_X1    g0357(.A(new_n542), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n264), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n540), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n297), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G190), .B(new_n540), .C1(new_n546), .C2(new_n264), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n550), .A2(KEYINPUT86), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT86), .B1(new_n550), .B2(new_n564), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(G20), .B1(new_n342), .B2(G97), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n476), .B1(G20), .B2(new_n541), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n288), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n288), .A3(KEYINPUT20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n291), .A2(new_n541), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT87), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n471), .B2(new_n541), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n505), .A2(KEYINPUT87), .A3(G116), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G303), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n264), .B1(new_n255), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n256), .A2(G257), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G264), .A2(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n545), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n486), .A2(new_n484), .ZN(new_n586));
  OAI211_X1 g0386(.A(G270), .B(new_n264), .C1(new_n482), .C2(new_n483), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n588), .A2(G169), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n579), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(KEYINPUT21), .A3(G169), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n585), .A2(new_n586), .A3(G179), .A4(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n590), .A2(new_n591), .B1(new_n594), .B2(new_n579), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n588), .A2(G200), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n379), .B2(new_n588), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n579), .B2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n230), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n599));
  NAND2_X1  g0399(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n545), .A2(new_n230), .A3(G87), .A4(new_n600), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT24), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT23), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n230), .B2(G107), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n459), .A2(KEYINPUT23), .A3(G20), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n542), .B2(new_n230), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n604), .B2(new_n609), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n288), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n291), .A2(new_n459), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT25), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(G107), .B2(new_n505), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G294), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n618), .C1(new_n479), .C2(G1698), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n265), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n485), .A2(G264), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n586), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n332), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n622), .A2(G179), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n620), .A2(new_n621), .A3(G190), .A4(new_n586), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(G200), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n612), .A2(new_n615), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n598), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n457), .A2(new_n502), .A3(new_n567), .A4(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n566), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n550), .A2(KEYINPUT86), .A3(new_n564), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n489), .ZN(new_n635));
  INV_X1    g0435(.A(new_n492), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n491), .B1(new_n481), .B2(new_n487), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n332), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n533), .A2(new_n534), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n549), .B1(new_n554), .B2(new_n563), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n635), .A2(new_n642), .A3(new_n638), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n549), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n628), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n595), .B2(new_n625), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n502), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n457), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n337), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n439), .A2(new_n441), .ZN(new_n653));
  INV_X1    g0453(.A(new_n436), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n333), .B(new_n319), .C1(new_n326), .C2(G179), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT89), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n331), .A2(new_n658), .A3(new_n333), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n449), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n445), .B1(new_n661), .B2(new_n447), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n422), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n406), .B(new_n410), .C1(new_n664), .C2(new_n400), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n652), .B1(new_n665), .B2(new_n304), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n651), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n289), .A2(new_n230), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n595), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT90), .Z(new_n675));
  OR2_X1    g0475(.A1(new_n625), .A2(new_n673), .ZN(new_n676));
  INV_X1    g0476(.A(new_n628), .ZN(new_n677));
  INV_X1    g0477(.A(new_n673), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n612), .B2(new_n615), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n625), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n676), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n579), .A2(new_n673), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n595), .B(new_n684), .C1(new_n579), .C2(new_n597), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n595), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n681), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(G399));
  NOR2_X1   g0490(.A1(new_n525), .A2(G116), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n233), .A2(new_n267), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n227), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n673), .B1(new_n640), .B2(new_n649), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n495), .A2(new_n496), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n501), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n625), .A2(new_n595), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n642), .A2(new_n628), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n639), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT92), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT92), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n648), .A2(new_n707), .A3(new_n639), .A4(new_n702), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n632), .A2(new_n643), .A3(new_n494), .A4(new_n633), .ZN(new_n709));
  INV_X1    g0509(.A(new_n645), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n494), .A2(new_n642), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT26), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n706), .A2(new_n708), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n698), .B1(new_n713), .B2(new_n678), .ZN(new_n714));
  INV_X1    g0514(.A(G330), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n636), .A2(new_n637), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n620), .A2(new_n621), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n593), .A3(new_n547), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n547), .A2(new_n330), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n488), .A2(new_n722), .A3(new_n588), .A4(new_n622), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT91), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n716), .A2(KEYINPUT30), .A3(new_n718), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n673), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n721), .A2(new_n725), .A3(new_n723), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n678), .A2(new_n728), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n567), .A2(new_n502), .A3(new_n630), .A4(new_n678), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n715), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n699), .A2(new_n714), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n696), .B1(new_n734), .B2(G1), .ZN(G364));
  XNOR2_X1  g0535(.A(new_n687), .B(KEYINPUT93), .ZN(new_n736));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n289), .B1(new_n738), .B2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n692), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n736), .B(new_n740), .C1(G330), .C2(new_n686), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT94), .ZN(new_n742));
  INV_X1    g0542(.A(new_n740), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n545), .A2(new_n233), .ZN(new_n744));
  INV_X1    g0544(.A(G355), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(G116), .B2(new_n233), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n228), .A2(new_n268), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n255), .A2(new_n233), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n248), .B2(G45), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n229), .B1(G20), .B2(new_n332), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n743), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n379), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n230), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n230), .A2(new_n330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n379), .ZN(new_n763));
  AOI22_X1  g0563(.A1(G294), .A2(new_n760), .B1(new_n763), .B2(G326), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT96), .Z(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n230), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n766), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(G311), .B1(new_n771), .B2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  INV_X1    g0573(.A(new_n761), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n774), .A2(new_n379), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n772), .B(new_n255), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n762), .A2(G190), .ZN(new_n778));
  XNOR2_X1  g0578(.A(KEYINPUT33), .B(G317), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT95), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n297), .A2(new_n769), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(new_n379), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n297), .A2(KEYINPUT95), .A3(G190), .A4(new_n769), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G303), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G283), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n765), .A2(new_n780), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n545), .B1(new_n209), .B2(new_n767), .C1(new_n776), .C2(new_n202), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G107), .B2(new_n788), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n759), .A2(new_n461), .ZN(new_n793));
  INV_X1    g0593(.A(new_n778), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n203), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n793), .B(new_n795), .C1(G50), .C2(new_n763), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n770), .A2(new_n353), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n792), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n785), .B1(new_n523), .B2(new_n524), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n790), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n757), .B1(new_n801), .B2(new_n754), .ZN(new_n802));
  INV_X1    g0602(.A(new_n753), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n686), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n742), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT97), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NAND4_X1  g0607(.A1(new_n657), .A2(new_n319), .A3(new_n659), .A4(new_n673), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n319), .A2(new_n673), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n334), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n697), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n334), .B2(new_n697), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n733), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n743), .B1(new_n813), .B2(new_n733), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(KEYINPUT98), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(KEYINPUT98), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n754), .A2(new_n751), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n743), .B1(new_n819), .B2(G77), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n794), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n793), .B(new_n822), .C1(G303), .C2(new_n763), .ZN(new_n823));
  INV_X1    g0623(.A(new_n788), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n307), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n255), .B1(new_n767), .B2(new_n541), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n776), .A2(new_n827), .B1(new_n770), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n823), .B(new_n830), .C1(new_n459), .C2(new_n785), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n775), .A2(G143), .B1(G159), .B2(new_n768), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(new_n763), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n834), .C1(new_n278), .C2(new_n794), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  NOR2_X1   g0636(.A1(new_n759), .A2(new_n202), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n255), .B(new_n837), .C1(G132), .C2(new_n771), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n824), .B2(new_n203), .C1(new_n785), .C2(new_n201), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n831), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n820), .B1(new_n840), .B2(new_n754), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n811), .B2(new_n752), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n817), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n738), .A2(new_n289), .ZN(new_n844));
  INV_X1    g0644(.A(new_n671), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n367), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n402), .B2(new_n384), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n367), .A2(KEYINPUT100), .A3(new_n408), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT100), .B1(new_n367), .B2(new_n408), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n846), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n340), .B1(new_n852), .B2(new_n366), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n408), .B2(new_n845), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n384), .B(new_n340), .C1(new_n361), .C2(new_n366), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n845), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(KEYINPUT38), .C1(new_n412), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT103), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n367), .A2(new_n408), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n846), .A3(new_n855), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n847), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n851), .A2(new_n865), .A3(KEYINPUT102), .ZN(new_n866));
  INV_X1    g0666(.A(new_n846), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n400), .B2(new_n411), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT102), .B1(new_n851), .B2(new_n865), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n861), .B(new_n862), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n851), .A2(new_n865), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n868), .A3(new_n866), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n861), .B1(new_n876), .B2(new_n862), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n860), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n727), .B(KEYINPUT31), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n732), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n451), .A2(new_n673), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n655), .B(new_n881), .C1(new_n662), .C2(new_n422), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n451), .B(new_n673), .C1(new_n450), .C2(new_n442), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(new_n811), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n880), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n412), .A2(new_n859), .ZN(new_n887));
  INV_X1    g0687(.A(new_n858), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n862), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n860), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n885), .A2(new_n890), .A3(new_n880), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n457), .A2(new_n880), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n715), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n656), .A2(new_n673), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n697), .B2(new_n334), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n882), .A2(new_n883), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n901), .A2(new_n890), .B1(new_n411), .B2(new_n671), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n860), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT103), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n906), .B2(new_n871), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n903), .B1(new_n889), .B2(new_n860), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n662), .A2(new_n422), .A3(new_n673), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n902), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n457), .B1(new_n714), .B2(new_n699), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n666), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n912), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n844), .B1(new_n897), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n897), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n227), .A2(G77), .A3(new_n357), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(G50), .B2(new_n203), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(G1), .A3(new_n737), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n465), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(G116), .A3(new_n231), .A4(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(KEYINPUT99), .B(KEYINPUT36), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n917), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT104), .ZN(G367));
  NOR2_X1   g0727(.A1(new_n554), .A2(new_n678), .ZN(new_n928));
  MUX2_X1   g0728(.A(new_n642), .B(new_n710), .S(new_n928), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT105), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n502), .B1(new_n495), .B2(new_n678), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n494), .A2(new_n673), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n682), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n639), .B1(new_n932), .B2(new_n625), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n678), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n689), .A2(new_n935), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n947));
  XNOR2_X1  g0747(.A(new_n692), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n683), .A2(new_n934), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT45), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n683), .A2(new_n934), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n688), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n675), .B(new_n681), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n687), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n736), .B2(new_n956), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n734), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n689), .A3(new_n953), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n949), .B1(new_n962), .B2(new_n734), .ZN(new_n963));
  INV_X1    g0763(.A(new_n739), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n946), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n244), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n755), .B1(new_n233), .B2(new_n315), .C1(new_n966), .C2(new_n748), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n743), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n768), .A2(G283), .B1(new_n771), .B2(G317), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n969), .B(new_n255), .C1(new_n580), .C2(new_n776), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G107), .A2(new_n760), .B1(new_n763), .B2(G311), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n827), .B2(new_n794), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(G97), .C2(new_n788), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n786), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n785), .B2(new_n541), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n759), .A2(new_n203), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n794), .A2(new_n353), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G143), .C2(new_n763), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n788), .A2(G77), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n255), .B1(new_n771), .B2(G137), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n775), .A2(G150), .B1(G50), .B2(new_n768), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n980), .B(new_n984), .C1(new_n202), .C2(new_n785), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT47), .Z(new_n987));
  INV_X1    g0787(.A(new_n754), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n968), .B1(new_n929), .B2(new_n803), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n965), .A2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n681), .A2(new_n753), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n691), .A2(new_n744), .B1(G107), .B2(new_n233), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n241), .A2(G45), .ZN(new_n993));
  INV_X1    g0793(.A(new_n691), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n994), .C1(G68), .C2(G77), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n281), .A2(G50), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n748), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n992), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n743), .B1(new_n1000), .B2(new_n756), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n508), .A2(new_n760), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n201), .B2(new_n776), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n786), .A2(G77), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n545), .B1(new_n770), .B2(new_n278), .C1(new_n203), .C2(new_n767), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n353), .A2(new_n834), .B1(new_n794), .B2(new_n281), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G97), .C2(new_n788), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n545), .B1(new_n771), .B2(G326), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n775), .A2(G317), .B1(G303), .B2(new_n768), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n828), .B2(new_n794), .C1(new_n773), .C2(new_n834), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n821), .B2(new_n759), .C1(new_n827), .C2(new_n785), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT49), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1010), .B1(new_n541), .B2(new_n824), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1001), .B1(new_n1018), .B2(new_n754), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n958), .A2(new_n964), .B1(new_n991), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n692), .B(KEYINPUT109), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n959), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n958), .A2(new_n734), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT110), .ZN(G393));
  NAND2_X1  g0825(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(new_n961), .Z(new_n1027));
  OAI211_X1 g0827(.A(new_n962), .B(new_n1021), .C1(new_n1027), .C2(new_n960), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n755), .B1(new_n461), .B2(new_n233), .C1(new_n251), .C2(new_n748), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G116), .A2(new_n760), .B1(new_n778), .B2(G303), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n255), .B1(new_n770), .B2(new_n773), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G294), .B2(new_n768), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(new_n459), .C2(new_n824), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n775), .A2(G311), .B1(new_n763), .B2(G317), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(G283), .C2(new_n786), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n255), .B(new_n825), .C1(G143), .C2(new_n771), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n217), .B2(new_n785), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT113), .Z(new_n1039));
  AOI22_X1  g0839(.A1(new_n775), .A2(G159), .B1(new_n763), .B2(G150), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n759), .A2(new_n209), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n305), .B2(new_n768), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n201), .B2(new_n794), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1042), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1036), .B1(new_n1039), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n743), .B(new_n1029), .C1(new_n1048), .C2(new_n988), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT114), .Z(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n753), .B2(new_n935), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1027), .B2(new_n964), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1028), .A2(new_n1052), .ZN(G390));
  AOI21_X1  g0853(.A(new_n715), .B1(new_n879), .B2(new_n732), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n885), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n643), .B1(new_n567), .B2(new_n494), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n646), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n705), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n334), .B(new_n678), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n898), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n910), .B1(new_n1062), .B2(new_n884), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n907), .A2(new_n1063), .A3(new_n908), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n860), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n906), .B2(new_n871), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n713), .A2(new_n811), .A3(new_n678), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n900), .B1(new_n1067), .B2(new_n1061), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1066), .A2(new_n910), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1056), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT115), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT115), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n1056), .C1(new_n1064), .C2(new_n1069), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n733), .A2(new_n811), .A3(new_n884), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n457), .A2(new_n1054), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n913), .A2(new_n666), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1054), .A2(new_n811), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n900), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1081), .A2(new_n1061), .A3(new_n1067), .A4(new_n1075), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n884), .B1(new_n733), .B2(new_n811), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1062), .B1(new_n1056), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1079), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1077), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1071), .A2(new_n1073), .A3(new_n1076), .A4(new_n1085), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1087), .A2(new_n1021), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n909), .A2(new_n751), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n771), .A2(G125), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n545), .B1(new_n824), .B2(new_n201), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT117), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT118), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G159), .A2(new_n760), .B1(new_n778), .B2(G137), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT54), .B(G143), .Z(new_n1099));
  AOI22_X1  g0899(.A1(new_n775), .A2(G132), .B1(new_n768), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1100), .C1(new_n1101), .C2(new_n834), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n786), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT53), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n785), .B2(new_n278), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1097), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n545), .B1(new_n771), .B2(G294), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n461), .B2(new_n767), .C1(new_n776), .C2(new_n541), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G68), .B2(new_n788), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n834), .A2(new_n821), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1043), .B(new_n1111), .C1(G107), .C2(new_n778), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(new_n307), .C2(new_n785), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n988), .B1(new_n1107), .B2(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n740), .B(new_n1114), .C1(new_n281), .C2(new_n818), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1091), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT119), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(KEYINPUT120), .C1(new_n739), .C2(new_n1077), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT116), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1087), .A2(new_n1120), .A3(new_n1021), .A4(new_n1088), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1077), .A2(new_n739), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n1117), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1090), .A2(new_n1119), .A3(new_n1121), .A4(new_n1124), .ZN(G378));
  NOR2_X1   g0925(.A1(G33), .A2(G41), .ZN(new_n1126));
  AOI211_X1 g0926(.A(G50), .B(new_n1126), .C1(new_n255), .C2(new_n267), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n794), .A2(new_n461), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n978), .B(new_n1128), .C1(G116), .C2(new_n763), .ZN(new_n1129));
  AOI211_X1 g0929(.A(G41), .B(new_n545), .C1(new_n771), .C2(G283), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n459), .B2(new_n776), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n508), .B2(new_n768), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n788), .A2(G58), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1129), .A2(new_n1132), .A3(new_n1005), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT58), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1135), .B2(new_n1134), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n776), .A2(new_n1101), .B1(new_n767), .B2(new_n833), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G132), .B2(new_n778), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n786), .A2(new_n1099), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(G150), .A2(new_n760), .B1(new_n763), .B2(G125), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n771), .A2(G124), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1126), .B(new_n1145), .C1(new_n824), .C2(new_n353), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n754), .B1(new_n1137), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n740), .B1(new_n201), .B2(new_n818), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n304), .A2(new_n337), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n295), .A2(new_n845), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT121), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT121), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1148), .B(new_n1149), .C1(new_n1161), .C2(new_n752), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n886), .A2(G330), .A3(new_n893), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1161), .A2(G330), .A3(new_n893), .A4(new_n886), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1165), .A2(new_n912), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n912), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1169), .B2(new_n964), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1021), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1079), .B(KEYINPUT122), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n1088), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT123), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT123), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1088), .A2(new_n1176), .A3(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1167), .A2(new_n1168), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1172), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1088), .A2(new_n1176), .A3(new_n1173), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1176), .B1(new_n1088), .B2(new_n1173), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1169), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1179), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1171), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1079), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1086), .A3(new_n948), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT124), .Z(new_n1192));
  OAI21_X1  g0992(.A(new_n743), .B1(new_n819), .B2(G68), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n778), .A2(new_n1099), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n201), .B2(new_n759), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G132), .B2(new_n763), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n255), .B1(new_n775), .B2(G137), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n768), .A2(G150), .B1(new_n771), .B2(G128), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1133), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(new_n353), .C2(new_n785), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n541), .A2(new_n794), .B1(new_n834), .B2(new_n827), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n255), .B1(new_n776), .B2(new_n821), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n767), .A2(new_n459), .B1(new_n770), .B2(new_n580), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n981), .A3(new_n1002), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n785), .A2(new_n461), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1193), .B1(new_n1207), .B2(new_n754), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n884), .B2(new_n752), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1189), .B2(new_n739), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1192), .A2(new_n1211), .ZN(G381));
  OR2_X1    g1012(.A1(G390), .A2(G387), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1124), .A2(new_n1089), .A3(new_n1119), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n1186), .A3(new_n1215), .A4(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n672), .A2(G213), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1186), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G407), .A2(G213), .A3(new_n1220), .ZN(G409));
  AOI21_X1  g1021(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1169), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1180), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1021), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G378), .B(new_n1170), .C1(new_n1222), .C2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1170), .B1(new_n1184), .B2(new_n949), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1216), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1190), .B2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1189), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1079), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1172), .B(new_n1085), .C1(new_n1190), .C2(new_n1230), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1211), .ZN(new_n1236));
  INV_X1    g1036(.A(G384), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(G384), .A3(new_n1211), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1228), .A2(new_n1218), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT62), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1219), .A2(G2897), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1238), .A2(new_n1239), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1186), .A2(G378), .B1(new_n1216), .B2(new_n1226), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1248), .B2(new_n1219), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT62), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1228), .A2(new_n1250), .A3(new_n1240), .A4(new_n1218), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1242), .A2(new_n1243), .A3(new_n1249), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G390), .A2(G387), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1213), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(G393), .B(new_n806), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1213), .A2(new_n1256), .A3(new_n1254), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1228), .A2(new_n1218), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1247), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT127), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1242), .A3(new_n1263), .A4(new_n1251), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1260), .A3(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1249), .B(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1241), .B(KEYINPUT63), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1243), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(G405));
  INV_X1    g1070(.A(new_n1216), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1225), .B1(new_n1186), .B2(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(new_n1240), .Z(new_n1273));
  XNOR2_X1  g1073(.A(new_n1267), .B(new_n1273), .ZN(G402));
endmodule


