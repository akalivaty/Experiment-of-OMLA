

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741;

  NOR2_X1 U372 ( .A1(n525), .A2(n385), .ZN(n529) );
  AND2_X1 U373 ( .A1(n368), .A2(n367), .ZN(n366) );
  OR2_X1 U374 ( .A1(n597), .A2(n474), .ZN(n367) );
  NOR2_X2 U375 ( .A1(n519), .A2(n520), .ZN(n540) );
  XNOR2_X2 U376 ( .A(n501), .B(n439), .ZN(n471) );
  NOR2_X1 U377 ( .A1(n386), .A2(n510), .ZN(n513) );
  XNOR2_X2 U378 ( .A(n361), .B(KEYINPUT19), .ZN(n574) );
  XNOR2_X2 U379 ( .A(n471), .B(n440), .ZN(n402) );
  XNOR2_X2 U380 ( .A(n711), .B(n421), .ZN(n697) );
  NOR2_X1 U381 ( .A1(n530), .A2(n661), .ZN(n531) );
  XNOR2_X2 U382 ( .A(n472), .B(n400), .ZN(n711) );
  NAND2_X1 U383 ( .A1(n533), .A2(n532), .ZN(n656) );
  INV_X1 U384 ( .A(KEYINPUT3), .ZN(n360) );
  XNOR2_X1 U385 ( .A(n384), .B(KEYINPUT35), .ZN(n733) );
  XNOR2_X1 U386 ( .A(n524), .B(KEYINPUT110), .ZN(n735) );
  NOR2_X2 U387 ( .A1(n536), .A2(n597), .ZN(n523) );
  XNOR2_X1 U388 ( .A(n380), .B(KEYINPUT39), .ZN(n596) );
  XNOR2_X1 U389 ( .A(n529), .B(n528), .ZN(n661) );
  XNOR2_X1 U390 ( .A(n521), .B(KEYINPUT6), .ZN(n546) );
  OR2_X1 U391 ( .A1(n628), .A2(G902), .ZN(n377) );
  XNOR2_X1 U392 ( .A(n401), .B(n445), .ZN(n400) );
  XNOR2_X1 U393 ( .A(n399), .B(n412), .ZN(n398) );
  XNOR2_X1 U394 ( .A(n360), .B(G113), .ZN(n399) );
  XNOR2_X1 U395 ( .A(n438), .B(n437), .ZN(n501) );
  XNOR2_X1 U396 ( .A(n413), .B(G104), .ZN(n445) );
  XNOR2_X1 U397 ( .A(n414), .B(KEYINPUT16), .ZN(n401) );
  XNOR2_X1 U398 ( .A(G146), .B(G125), .ZN(n447) );
  XNOR2_X1 U399 ( .A(G131), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U400 ( .A(G101), .B(G119), .ZN(n412) );
  XNOR2_X2 U401 ( .A(n352), .B(n353), .ZN(n559) );
  NOR2_X1 U402 ( .A1(n702), .A2(G902), .ZN(n352) );
  XOR2_X1 U403 ( .A(KEYINPUT68), .B(G469), .Z(n353) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n484) );
  XNOR2_X1 U405 ( .A(G140), .B(G137), .ZN(n449) );
  INV_X1 U406 ( .A(G134), .ZN(n437) );
  AND2_X1 U407 ( .A1(n735), .A2(n383), .ZN(n381) );
  INV_X1 U408 ( .A(KEYINPUT15), .ZN(n422) );
  NOR2_X1 U409 ( .A1(G237), .A2(G902), .ZN(n410) );
  XNOR2_X1 U410 ( .A(G137), .B(G146), .ZN(n466) );
  NOR2_X1 U411 ( .A1(n374), .A2(G953), .ZN(n453) );
  XOR2_X1 U412 ( .A(G131), .B(G140), .Z(n486) );
  XNOR2_X1 U413 ( .A(G113), .B(G143), .ZN(n479) );
  NAND2_X1 U414 ( .A1(n476), .A2(n597), .ZN(n385) );
  NAND2_X1 U415 ( .A1(n406), .A2(KEYINPUT100), .ZN(n368) );
  NAND2_X1 U416 ( .A1(n375), .A2(G953), .ZN(n548) );
  INV_X1 U417 ( .A(n547), .ZN(n375) );
  BUF_X1 U418 ( .A(n521), .Z(n670) );
  XNOR2_X1 U419 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n448) );
  XNOR2_X1 U420 ( .A(G119), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U421 ( .A(G128), .B(G110), .ZN(n452) );
  NOR2_X1 U422 ( .A1(n535), .A2(n668), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n511), .B(KEYINPUT22), .ZN(n512) );
  XNOR2_X1 U424 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U425 ( .A(n405), .B(n617), .ZN(n404) );
  NOR2_X1 U426 ( .A1(n627), .A2(n490), .ZN(n405) );
  AND2_X1 U427 ( .A1(n393), .A2(n391), .ZN(n390) );
  NOR2_X1 U428 ( .A1(n392), .A2(n710), .ZN(n391) );
  XNOR2_X1 U429 ( .A(n595), .B(n594), .ZN(n379) );
  NOR2_X1 U430 ( .A1(n592), .A2(n591), .ZN(n595) );
  XOR2_X1 U431 ( .A(KEYINPUT4), .B(KEYINPUT18), .Z(n415) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n428) );
  XNOR2_X1 U433 ( .A(n425), .B(n424), .ZN(n426) );
  INV_X1 U434 ( .A(G902), .ZN(n503) );
  XNOR2_X1 U435 ( .A(n362), .B(n471), .ZN(n621) );
  XNOR2_X1 U436 ( .A(n472), .B(n470), .ZN(n362) );
  AND2_X1 U437 ( .A1(n379), .A2(n603), .ZN(n725) );
  XNOR2_X1 U438 ( .A(n489), .B(n488), .ZN(n616) );
  AND2_X1 U439 ( .A1(n551), .A2(n408), .ZN(n552) );
  AND2_X1 U440 ( .A1(n546), .A2(n664), .ZN(n551) );
  NAND2_X1 U441 ( .A1(n407), .A2(n365), .ZN(n364) );
  NOR2_X1 U442 ( .A1(n558), .A2(n557), .ZN(n561) );
  XNOR2_X1 U443 ( .A(n521), .B(KEYINPUT109), .ZN(n568) );
  INV_X1 U444 ( .A(G953), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n456), .B(n457), .ZN(n628) );
  XNOR2_X1 U446 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U447 ( .A(n402), .B(n446), .ZN(n702) );
  XNOR2_X1 U448 ( .A(G146), .B(KEYINPUT75), .ZN(n442) );
  AND2_X1 U449 ( .A1(n596), .A2(n583), .ZN(n585) );
  XNOR2_X1 U450 ( .A(n369), .B(KEYINPUT32), .ZN(n739) );
  NOR2_X1 U451 ( .A1(n536), .A2(n370), .ZN(n369) );
  INV_X1 U452 ( .A(KEYINPUT76), .ZN(n371) );
  NAND2_X1 U453 ( .A1(n404), .A2(n396), .ZN(n403) );
  INV_X1 U454 ( .A(KEYINPUT56), .ZN(n394) );
  XOR2_X1 U455 ( .A(G122), .B(G104), .Z(n354) );
  AND2_X1 U456 ( .A1(n569), .A2(n465), .ZN(n476) );
  XOR2_X1 U457 ( .A(n600), .B(n581), .Z(n355) );
  AND2_X1 U458 ( .A1(n560), .A2(n355), .ZN(n356) );
  AND2_X1 U459 ( .A1(n603), .A2(KEYINPUT2), .ZN(n357) );
  INV_X1 U460 ( .A(G234), .ZN(n374) );
  INV_X1 U461 ( .A(KEYINPUT100), .ZN(n474) );
  AND2_X1 U462 ( .A1(n397), .A2(G210), .ZN(n358) );
  INV_X1 U463 ( .A(n699), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n697), .B(n698), .ZN(n699) );
  XOR2_X1 U465 ( .A(KEYINPUT66), .B(KEYINPUT60), .Z(n359) );
  INV_X1 U466 ( .A(n710), .ZN(n396) );
  XNOR2_X2 U467 ( .A(n398), .B(n411), .ZN(n472) );
  NAND2_X1 U468 ( .A1(n545), .A2(n653), .ZN(n361) );
  XNOR2_X1 U469 ( .A(n513), .B(n512), .ZN(n536) );
  INV_X1 U470 ( .A(n733), .ZN(n382) );
  XNOR2_X2 U471 ( .A(n363), .B(KEYINPUT31), .ZN(n646) );
  NOR2_X2 U472 ( .A1(n675), .A2(n386), .ZN(n363) );
  XNOR2_X1 U473 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X2 U474 ( .A(n505), .B(n504), .ZN(n533) );
  INV_X1 U475 ( .A(n597), .ZN(n668) );
  NAND2_X1 U476 ( .A1(n366), .A2(n364), .ZN(n675) );
  AND2_X1 U477 ( .A1(n597), .A2(n474), .ZN(n365) );
  XNOR2_X2 U478 ( .A(n559), .B(KEYINPUT1), .ZN(n597) );
  XNOR2_X1 U479 ( .A(n372), .B(n371), .ZN(n370) );
  NAND2_X1 U480 ( .A1(n373), .A2(n506), .ZN(n507) );
  NAND2_X1 U481 ( .A1(n646), .A2(n633), .ZN(n373) );
  NAND2_X1 U482 ( .A1(n376), .A2(G227), .ZN(n441) );
  NAND2_X1 U483 ( .A1(n376), .A2(G224), .ZN(n419) );
  NAND2_X1 U484 ( .A1(n726), .A2(n376), .ZN(n732) );
  XNOR2_X2 U485 ( .A(n377), .B(n462), .ZN(n569) );
  NAND2_X1 U486 ( .A1(n379), .A2(n357), .ZN(n378) );
  XNOR2_X1 U487 ( .A(n378), .B(KEYINPUT85), .ZN(n610) );
  NAND2_X1 U488 ( .A1(n561), .A2(n560), .ZN(n582) );
  NAND2_X1 U489 ( .A1(n561), .A2(n356), .ZN(n380) );
  NAND2_X1 U490 ( .A1(n382), .A2(n381), .ZN(n538) );
  INV_X1 U491 ( .A(n739), .ZN(n383) );
  NAND2_X1 U492 ( .A1(n387), .A2(n563), .ZN(n384) );
  NOR2_X2 U493 ( .A1(n624), .A2(n710), .ZN(n626) );
  XNOR2_X1 U494 ( .A(n403), .B(n359), .ZN(G60) );
  XNOR2_X1 U495 ( .A(n386), .B(n475), .ZN(n530) );
  XNOR2_X2 U496 ( .A(n436), .B(KEYINPUT0), .ZN(n386) );
  XNOR2_X1 U497 ( .A(n531), .B(KEYINPUT34), .ZN(n387) );
  NAND2_X1 U498 ( .A1(n696), .A2(n358), .ZN(n393) );
  NAND2_X1 U499 ( .A1(n390), .A2(n388), .ZN(n395) );
  NAND2_X1 U500 ( .A1(n389), .A2(n699), .ZN(n388) );
  INV_X1 U501 ( .A(n696), .ZN(n389) );
  NOR2_X1 U502 ( .A1(n397), .A2(G210), .ZN(n392) );
  XNOR2_X1 U503 ( .A(n395), .B(n394), .ZN(G51) );
  XNOR2_X1 U504 ( .A(n402), .B(n724), .ZN(n727) );
  NOR2_X2 U505 ( .A1(n667), .A2(n670), .ZN(n407) );
  INV_X1 U506 ( .A(n407), .ZN(n406) );
  BUF_X1 U507 ( .A(n609), .Z(n714) );
  XNOR2_X1 U508 ( .A(n542), .B(n541), .ZN(n609) );
  XNOR2_X1 U509 ( .A(n427), .B(n426), .ZN(n545) );
  AND2_X1 U510 ( .A1(n567), .A2(n653), .ZN(n408) );
  INV_X1 U511 ( .A(KEYINPUT108), .ZN(n517) );
  INV_X1 U512 ( .A(KEYINPUT17), .ZN(n416) );
  INV_X1 U513 ( .A(KEYINPUT9), .ZN(n497) );
  XNOR2_X1 U514 ( .A(n593), .B(KEYINPUT48), .ZN(n594) );
  XNOR2_X1 U515 ( .A(n487), .B(n724), .ZN(n488) );
  INV_X1 U516 ( .A(KEYINPUT79), .ZN(n424) );
  INV_X1 U517 ( .A(KEYINPUT38), .ZN(n581) );
  INV_X1 U518 ( .A(G475), .ZN(n490) );
  INV_X1 U519 ( .A(KEYINPUT41), .ZN(n586) );
  XNOR2_X1 U520 ( .A(n587), .B(n586), .ZN(n651) );
  XNOR2_X1 U521 ( .A(n493), .B(n492), .ZN(n508) );
  INV_X1 U522 ( .A(G952), .ZN(n409) );
  AND2_X1 U523 ( .A1(n409), .A2(G953), .ZN(n710) );
  AND2_X1 U524 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n520) );
  XOR2_X1 U525 ( .A(KEYINPUT74), .B(n410), .Z(n423) );
  NAND2_X1 U526 ( .A1(n423), .A2(G214), .ZN(n653) );
  XNOR2_X1 U527 ( .A(G116), .B(KEYINPUT69), .ZN(n411) );
  XOR2_X1 U528 ( .A(KEYINPUT73), .B(G122), .Z(n414) );
  XNOR2_X1 U529 ( .A(G110), .B(G107), .ZN(n413) );
  XNOR2_X1 U530 ( .A(n447), .B(n415), .ZN(n418) );
  XNOR2_X2 U531 ( .A(G143), .B(G128), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n438), .B(n416), .ZN(n417) );
  XNOR2_X1 U533 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U534 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U535 ( .A(n422), .B(G902), .ZN(n605) );
  NOR2_X1 U536 ( .A1(n697), .A2(n605), .ZN(n427) );
  NAND2_X1 U537 ( .A1(G210), .A2(n423), .ZN(n425) );
  XNOR2_X1 U538 ( .A(n428), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U539 ( .A(KEYINPUT14), .B(n429), .ZN(n431) );
  NAND2_X1 U540 ( .A1(n431), .A2(G952), .ZN(n430) );
  XOR2_X1 U541 ( .A(KEYINPUT91), .B(n430), .Z(n683) );
  NOR2_X1 U542 ( .A1(G953), .A2(n683), .ZN(n550) );
  NAND2_X1 U543 ( .A1(n431), .A2(G902), .ZN(n432) );
  XNOR2_X1 U544 ( .A(KEYINPUT94), .B(n432), .ZN(n547) );
  XOR2_X1 U545 ( .A(G898), .B(KEYINPUT92), .Z(n719) );
  NAND2_X1 U546 ( .A1(n719), .A2(G953), .ZN(n433) );
  XOR2_X1 U547 ( .A(KEYINPUT93), .B(n433), .Z(n713) );
  NOR2_X1 U548 ( .A1(n547), .A2(n713), .ZN(n434) );
  OR2_X1 U549 ( .A1(n550), .A2(n434), .ZN(n435) );
  NAND2_X1 U550 ( .A1(n574), .A2(n435), .ZN(n436) );
  INV_X1 U551 ( .A(n449), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n441), .B(G101), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U554 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U555 ( .A(n447), .B(KEYINPUT10), .ZN(n724) );
  XNOR2_X1 U556 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U557 ( .A(n724), .B(n450), .ZN(n457) );
  XNOR2_X1 U558 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U559 ( .A(n453), .B(KEYINPUT8), .ZN(n494) );
  NAND2_X1 U560 ( .A1(n494), .A2(G221), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n455), .B(n454), .ZN(n456) );
  OR2_X1 U562 ( .A1(n605), .A2(n374), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n458), .B(KEYINPUT20), .ZN(n463) );
  NAND2_X1 U564 ( .A1(n463), .A2(G217), .ZN(n461) );
  XNOR2_X1 U565 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n463), .A2(G221), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n464), .B(KEYINPUT21), .ZN(n663) );
  INV_X1 U570 ( .A(n663), .ZN(n465) );
  INV_X1 U571 ( .A(n476), .ZN(n667) );
  XOR2_X1 U572 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n467) );
  XNOR2_X1 U573 ( .A(n467), .B(n466), .ZN(n469) );
  NAND2_X1 U574 ( .A1(n484), .A2(G210), .ZN(n468) );
  XNOR2_X1 U575 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U576 ( .A1(n621), .A2(n503), .ZN(n473) );
  INV_X1 U577 ( .A(G472), .ZN(n620) );
  XNOR2_X2 U578 ( .A(n473), .B(n620), .ZN(n521) );
  INV_X1 U579 ( .A(KEYINPUT95), .ZN(n475) );
  AND2_X1 U580 ( .A1(n670), .A2(n476), .ZN(n477) );
  NAND2_X1 U581 ( .A1(n477), .A2(n559), .ZN(n478) );
  OR2_X1 U582 ( .A1(n530), .A2(n478), .ZN(n633) );
  XNOR2_X1 U583 ( .A(n354), .B(n479), .ZN(n483) );
  XOR2_X1 U584 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n481) );
  XNOR2_X1 U585 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U587 ( .A(n483), .B(n482), .Z(n489) );
  NAND2_X1 U588 ( .A1(G214), .A2(n484), .ZN(n485) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U590 ( .A1(n616), .A2(G902), .ZN(n493) );
  XNOR2_X1 U591 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n491) );
  XOR2_X1 U592 ( .A(G107), .B(KEYINPUT7), .Z(n496) );
  NAND2_X1 U593 ( .A1(n494), .A2(G217), .ZN(n495) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U595 ( .A(G116), .B(G122), .ZN(n498) );
  XNOR2_X1 U596 ( .A(n501), .B(n502), .ZN(n706) );
  NAND2_X1 U597 ( .A1(n706), .A2(n503), .ZN(n505) );
  XOR2_X1 U598 ( .A(KEYINPUT104), .B(G478), .Z(n504) );
  NOR2_X1 U599 ( .A1(n508), .A2(n533), .ZN(n644) );
  AND2_X1 U600 ( .A1(n508), .A2(n533), .ZN(n583) );
  NOR2_X1 U601 ( .A1(n644), .A2(n583), .ZN(n658) );
  INV_X1 U602 ( .A(n658), .ZN(n506) );
  XNOR2_X1 U603 ( .A(n507), .B(KEYINPUT105), .ZN(n516) );
  INV_X1 U604 ( .A(n508), .ZN(n532) );
  NOR2_X1 U605 ( .A1(n663), .A2(n656), .ZN(n509) );
  XOR2_X1 U606 ( .A(KEYINPUT106), .B(n509), .Z(n510) );
  XNOR2_X1 U607 ( .A(KEYINPUT65), .B(KEYINPUT72), .ZN(n511) );
  INV_X1 U608 ( .A(n569), .ZN(n664) );
  NOR2_X1 U609 ( .A1(n546), .A2(n664), .ZN(n514) );
  NAND2_X1 U610 ( .A1(n523), .A2(n514), .ZN(n515) );
  XNOR2_X1 U611 ( .A(n515), .B(KEYINPUT107), .ZN(n734) );
  NOR2_X1 U612 ( .A1(n516), .A2(n734), .ZN(n518) );
  XNOR2_X1 U613 ( .A(n518), .B(n517), .ZN(n519) );
  NOR2_X1 U614 ( .A1(n568), .A2(n569), .ZN(n522) );
  NAND2_X1 U615 ( .A1(n523), .A2(n522), .ZN(n524) );
  INV_X1 U616 ( .A(n546), .ZN(n525) );
  XOR2_X1 U617 ( .A(KEYINPUT88), .B(KEYINPUT70), .Z(n527) );
  XNOR2_X1 U618 ( .A(KEYINPUT111), .B(KEYINPUT33), .ZN(n526) );
  XNOR2_X1 U619 ( .A(n527), .B(n526), .ZN(n528) );
  NOR2_X1 U620 ( .A1(n533), .A2(n532), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT77), .B(n546), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n534), .A2(n664), .ZN(n535) );
  NOR2_X1 U623 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U624 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U625 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U626 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n541) );
  NAND2_X1 U627 ( .A1(n609), .A2(n605), .ZN(n544) );
  INV_X1 U628 ( .A(KEYINPUT82), .ZN(n543) );
  XNOR2_X1 U629 ( .A(n544), .B(n543), .ZN(n604) );
  INV_X1 U630 ( .A(n545), .ZN(n600) );
  XNOR2_X1 U631 ( .A(n583), .B(KEYINPUT112), .ZN(n632) );
  INV_X1 U632 ( .A(n632), .ZN(n618) );
  NOR2_X1 U633 ( .A1(G900), .A2(n548), .ZN(n549) );
  NOR2_X1 U634 ( .A1(n550), .A2(n549), .ZN(n558) );
  NOR2_X1 U635 ( .A1(n663), .A2(n558), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n632), .A2(n552), .ZN(n598) );
  NOR2_X1 U637 ( .A1(n600), .A2(n598), .ZN(n553) );
  XOR2_X1 U638 ( .A(KEYINPUT36), .B(n553), .Z(n554) );
  NOR2_X1 U639 ( .A1(n554), .A2(n668), .ZN(n555) );
  XNOR2_X1 U640 ( .A(n555), .B(KEYINPUT114), .ZN(n737) );
  NAND2_X1 U641 ( .A1(n658), .A2(KEYINPUT47), .ZN(n564) );
  NAND2_X1 U642 ( .A1(n568), .A2(n653), .ZN(n556) );
  XNOR2_X1 U643 ( .A(n556), .B(KEYINPUT30), .ZN(n557) );
  INV_X1 U644 ( .A(n559), .ZN(n572) );
  NOR2_X1 U645 ( .A1(n572), .A2(n667), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n600), .A2(n582), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n641) );
  NAND2_X1 U648 ( .A1(n564), .A2(n641), .ZN(n565) );
  XNOR2_X1 U649 ( .A(KEYINPUT80), .B(n565), .ZN(n566) );
  NOR2_X1 U650 ( .A1(n737), .A2(n566), .ZN(n580) );
  INV_X1 U651 ( .A(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n570) );
  NOR2_X1 U653 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U654 ( .A(KEYINPUT28), .B(n571), .Z(n573) );
  NOR2_X1 U655 ( .A1(n573), .A2(n572), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n588), .A2(n574), .ZN(n575) );
  XOR2_X1 U657 ( .A(KEYINPUT78), .B(n575), .Z(n642) );
  XNOR2_X1 U658 ( .A(n576), .B(n642), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n576), .A2(n658), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n592) );
  XNOR2_X1 U662 ( .A(KEYINPUT40), .B(KEYINPUT113), .ZN(n584) );
  XNOR2_X1 U663 ( .A(n585), .B(n584), .ZN(n740) );
  NAND2_X1 U664 ( .A1(n355), .A2(n653), .ZN(n657) );
  NOR2_X1 U665 ( .A1(n656), .A2(n657), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n651), .A2(n588), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n589), .B(KEYINPUT42), .ZN(n741) );
  NAND2_X1 U668 ( .A1(n740), .A2(n741), .ZN(n590) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT46), .ZN(n591) );
  XOR2_X1 U670 ( .A(KEYINPUT86), .B(KEYINPUT67), .Z(n593) );
  NAND2_X1 U671 ( .A1(n596), .A2(n644), .ZN(n649) );
  OR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT43), .ZN(n601) );
  AND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n650) );
  INV_X1 U675 ( .A(n650), .ZN(n602) );
  AND2_X1 U676 ( .A1(n649), .A2(n602), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n725), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT83), .B(n605), .Z(n606) );
  NAND2_X1 U679 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n714), .A2(n610), .ZN(n684) );
  NAND2_X1 U682 ( .A1(n611), .A2(n684), .ZN(n612) );
  XNOR2_X2 U683 ( .A(n612), .B(KEYINPUT64), .ZN(n627) );
  XOR2_X1 U684 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n614) );
  XNOR2_X1 U685 ( .A(KEYINPUT122), .B(KEYINPUT89), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X1 U688 ( .A1(n646), .A2(n618), .ZN(n619) );
  XOR2_X1 U689 ( .A(G113), .B(n619), .Z(G15) );
  NOR2_X1 U690 ( .A1(n627), .A2(n620), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n621), .B(KEYINPUT62), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U693 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(G57) );
  INV_X2 U695 ( .A(n627), .ZN(n696) );
  NAND2_X1 U696 ( .A1(n696), .A2(G217), .ZN(n630) );
  XNOR2_X1 U697 ( .A(n628), .B(KEYINPUT124), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n631), .A2(n710), .ZN(G66) );
  INV_X1 U700 ( .A(n633), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n632), .A2(n635), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(G104), .ZN(G6) );
  XOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  NAND2_X1 U704 ( .A1(n635), .A2(n644), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(G107), .B(n638), .ZN(G9) );
  XOR2_X1 U707 ( .A(G128), .B(KEYINPUT29), .Z(n640) );
  NAND2_X1 U708 ( .A1(n644), .A2(n642), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(G30) );
  XNOR2_X1 U710 ( .A(G143), .B(n641), .ZN(G45) );
  NAND2_X1 U711 ( .A1(n632), .A2(n642), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(G146), .ZN(G48) );
  INV_X1 U713 ( .A(n644), .ZN(n645) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT116), .B(n647), .Z(n648) );
  XNOR2_X1 U716 ( .A(G116), .B(n648), .ZN(G18) );
  XNOR2_X1 U717 ( .A(G134), .B(n649), .ZN(G36) );
  XOR2_X1 U718 ( .A(G140), .B(n650), .Z(G42) );
  INV_X1 U719 ( .A(n651), .ZN(n678) );
  NOR2_X1 U720 ( .A1(n661), .A2(n678), .ZN(n652) );
  NOR2_X1 U721 ( .A1(G953), .A2(n652), .ZN(n693) );
  NOR2_X1 U722 ( .A1(n355), .A2(n653), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n654), .B(KEYINPUT118), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n680) );
  NAND2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U729 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n665) );
  XNOR2_X1 U730 ( .A(n666), .B(n665), .ZN(n673) );
  NAND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U732 ( .A(KEYINPUT50), .B(n669), .ZN(n671) );
  NAND2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U735 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U736 ( .A(n676), .B(KEYINPUT51), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U738 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U739 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U740 ( .A1(n683), .A2(n682), .ZN(n691) );
  INV_X1 U741 ( .A(n684), .ZN(n689) );
  OR2_X1 U742 ( .A1(n714), .A2(KEYINPUT2), .ZN(n687) );
  NOR2_X1 U743 ( .A1(n725), .A2(KEYINPUT2), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT81), .ZN(n686) );
  NAND2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U749 ( .A(n694), .B(KEYINPUT119), .ZN(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT53), .B(n695), .ZN(G75) );
  XOR2_X1 U751 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n698) );
  NAND2_X1 U752 ( .A1(n696), .A2(G469), .ZN(n704) );
  XOR2_X1 U753 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XNOR2_X1 U754 ( .A(n700), .B(KEYINPUT120), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U757 ( .A1(n710), .A2(n705), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n696), .A2(G478), .ZN(n708) );
  XNOR2_X1 U759 ( .A(n706), .B(KEYINPUT123), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U761 ( .A1(n710), .A2(n709), .ZN(G63) );
  XOR2_X1 U762 ( .A(KEYINPUT126), .B(n711), .Z(n712) );
  NAND2_X1 U763 ( .A1(n713), .A2(n712), .ZN(n723) );
  INV_X1 U764 ( .A(n714), .ZN(n715) );
  NOR2_X1 U765 ( .A1(n715), .A2(G953), .ZN(n721) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n716) );
  XNOR2_X1 U767 ( .A(n716), .B(KEYINPUT61), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n717), .B(KEYINPUT125), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U770 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n725), .B(n727), .ZN(n726) );
  XOR2_X1 U773 ( .A(G227), .B(n727), .Z(n728) );
  NAND2_X1 U774 ( .A1(n728), .A2(G900), .ZN(n729) );
  XOR2_X1 U775 ( .A(KEYINPUT127), .B(n729), .Z(n730) );
  NAND2_X1 U776 ( .A1(G953), .A2(n730), .ZN(n731) );
  NAND2_X1 U777 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U778 ( .A(n733), .B(G122), .Z(G24) );
  XOR2_X1 U779 ( .A(G101), .B(n734), .Z(G3) );
  XOR2_X1 U780 ( .A(G110), .B(n735), .Z(n736) );
  XNOR2_X1 U781 ( .A(KEYINPUT115), .B(n736), .ZN(G12) );
  XNOR2_X1 U782 ( .A(G125), .B(KEYINPUT37), .ZN(n738) );
  XNOR2_X1 U783 ( .A(n738), .B(n737), .ZN(G27) );
  XOR2_X1 U784 ( .A(G119), .B(n739), .Z(G21) );
  XNOR2_X1 U785 ( .A(n740), .B(G131), .ZN(G33) );
  XNOR2_X1 U786 ( .A(G137), .B(n741), .ZN(G39) );
endmodule

