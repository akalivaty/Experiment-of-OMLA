//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G58), .A2(G232), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n217), .A2(new_n227), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G68), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n213), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT70), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n218), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n248), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT11), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n247), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n205), .A2(G20), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n259), .A2(G68), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT12), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  AND4_X1   g0065(.A1(KEYINPUT12), .A2(new_n218), .A3(G20), .A4(new_n265), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n261), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n255), .A2(KEYINPUT11), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT71), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n256), .A2(new_n267), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT71), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n272), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  OAI211_X1 g0076(.A(G1), .B(G13), .C1(new_n252), .C2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G232), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G1698), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n280), .B(new_n282), .C1(G226), .C2(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G97), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT67), .A2(G41), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT67), .A2(G41), .ZN(new_n290));
  NOR3_X1   g0090(.A1(new_n289), .A2(new_n290), .A3(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n205), .A2(G274), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n219), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT13), .B1(new_n285), .B2(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(G169), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n298), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(new_n298), .B2(G169), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n275), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n268), .A2(new_n270), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G200), .ZN(new_n309));
  INV_X1    g0109(.A(new_n298), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n259), .A2(G50), .A3(new_n260), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G50), .B2(new_n257), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT8), .B(G58), .Z(new_n317));
  AOI22_X1  g0117(.A1(new_n317), .A2(new_n253), .B1(G150), .B2(new_n249), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n248), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT9), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n291), .A2(new_n292), .ZN(new_n324));
  INV_X1    g0124(.A(new_n288), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n325), .A2(G226), .ZN(new_n326));
  AOI21_X1  g0126(.A(G1698), .B1(new_n278), .B2(new_n279), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n327), .A2(G222), .B1(new_n330), .B2(G77), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n280), .A2(G1698), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT68), .B(G223), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n277), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n324), .B(new_n326), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G190), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n309), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n323), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT10), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n323), .A2(new_n341), .A3(new_n337), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n336), .A2(new_n301), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n322), .B1(new_n336), .B2(G169), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n317), .B(KEYINPUT69), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n249), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  INV_X1    g0149(.A(new_n253), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n348), .B1(new_n206), .B2(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n247), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n259), .A2(G77), .A3(new_n260), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G77), .B2(new_n257), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n324), .B1(G244), .B2(new_n325), .ZN(new_n358));
  INV_X1    g0158(.A(G107), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n332), .A2(new_n219), .B1(new_n359), .B2(new_n280), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(G232), .B2(new_n327), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n358), .B1(new_n361), .B2(new_n277), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(G179), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n362), .A2(new_n305), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(G200), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n367), .A2(new_n353), .A3(new_n356), .A4(new_n368), .ZN(new_n369));
  AND4_X1   g0169(.A1(new_n343), .A2(new_n346), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n259), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n317), .A2(new_n260), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(new_n257), .B2(new_n317), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  INV_X1    g0175(.A(G58), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n202), .B1(new_n218), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n278), .A2(new_n206), .A3(new_n279), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n279), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n218), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT74), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT74), .B(new_n218), .C1(new_n381), .C2(new_n382), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n375), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n330), .A2(new_n380), .A3(new_n206), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n379), .A2(KEYINPUT7), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G68), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n377), .A2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n249), .A2(G159), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT16), .A4(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n393), .A2(new_n247), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n387), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n387), .B2(new_n394), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n374), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n288), .A2(new_n281), .B1(new_n291), .B2(new_n292), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  OR2_X1    g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  INV_X1    g0201(.A(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(G226), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G87), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n403), .A2(new_n330), .B1(new_n252), .B2(new_n404), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n399), .A2(new_n400), .B1(new_n405), .B2(new_n335), .ZN(new_n406));
  OAI221_X1 g0206(.A(KEYINPUT76), .B1(new_n291), .B2(new_n292), .C1(new_n288), .C2(new_n281), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G179), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n364), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n398), .A2(new_n413), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT78), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n399), .A2(new_n400), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n335), .ZN(new_n419));
  AND4_X1   g0219(.A1(new_n305), .A2(new_n418), .A3(new_n407), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(G200), .B1(new_n406), .B2(new_n407), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT65), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G68), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n201), .B1(new_n426), .B2(G58), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n392), .B1(new_n427), .B2(new_n206), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n328), .A2(new_n329), .A3(G20), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT7), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT73), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n382), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n426), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n428), .B1(KEYINPUT74), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n386), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT16), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n393), .A2(new_n247), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT75), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n387), .A2(new_n394), .A3(new_n395), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n373), .B(new_n422), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n417), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n420), .A2(new_n421), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n374), .B(new_n446), .C1(new_n396), .C2(new_n397), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n447), .A2(KEYINPUT78), .A3(KEYINPUT17), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n447), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT77), .B1(new_n447), .B2(KEYINPUT17), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n445), .A2(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n314), .A2(new_n370), .A3(new_n416), .A4(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT79), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n289), .B2(new_n290), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n205), .A2(G45), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n455), .A2(KEYINPUT85), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT85), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT86), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT85), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n276), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT67), .A2(G41), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT5), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(new_n456), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT86), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n455), .A2(KEYINPUT85), .A3(new_n457), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n277), .B(G274), .C1(new_n454), .C2(G41), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n460), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G179), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n466), .A2(new_n468), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n454), .A2(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(new_n277), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G250), .B(new_n402), .C1(new_n328), .C2(new_n329), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT95), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n252), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n335), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT96), .B1(new_n473), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n470), .B1(new_n474), .B2(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n301), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT96), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n487), .A2(new_n488), .A3(new_n476), .A4(new_n483), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n472), .A2(new_n476), .A3(new_n483), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G169), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n485), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT97), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT97), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n485), .A2(new_n489), .A3(new_n494), .A4(new_n491), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n206), .B2(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n359), .A2(KEYINPUT23), .A3(G20), .ZN(new_n498));
  AND2_X1   g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n498), .B1(new_n206), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(KEYINPUT93), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT93), .B1(new_n501), .B2(KEYINPUT92), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n206), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(G20), .B1(new_n278), .B2(new_n279), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n503), .B1(new_n507), .B2(G87), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT94), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n505), .B(KEYINPUT93), .C1(KEYINPUT92), .C2(new_n501), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n507), .A2(G87), .A3(new_n503), .A4(new_n502), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT94), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n500), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n509), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n509), .B2(new_n513), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n247), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n205), .A2(G33), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n257), .A2(new_n518), .A3(new_n213), .A4(new_n246), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(G107), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n257), .A2(G107), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT25), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n493), .A2(new_n495), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT98), .ZN(new_n527));
  INV_X1    g0327(.A(new_n525), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n490), .A2(new_n309), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n472), .A2(new_n476), .A3(new_n483), .A4(new_n305), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n527), .B1(new_n526), .B2(new_n532), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT87), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n280), .A2(G244), .A3(new_n402), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  XOR2_X1   g0340(.A(new_n540), .B(KEYINPUT84), .Z(new_n541));
  NAND3_X1  g0341(.A1(new_n327), .A2(KEYINPUT4), .A3(G244), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n539), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n486), .A2(new_n469), .B1(new_n335), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n277), .C1(new_n474), .C2(new_n475), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n536), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n541), .A3(new_n543), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT4), .B1(new_n327), .B2(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n335), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n472), .A2(new_n546), .A3(new_n536), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n364), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n472), .A2(new_n546), .A3(new_n550), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(G179), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(G97), .B(G107), .ZN(new_n557));
  OR2_X1    g0357(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT80), .A2(KEYINPUT6), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n359), .A2(G97), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(KEYINPUT81), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(KEYINPUT81), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(G20), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n435), .A2(G107), .B1(G77), .B2(new_n249), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n248), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n258), .A2(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n520), .A2(new_n521), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(G97), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n553), .A2(new_n556), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n554), .A2(KEYINPUT87), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(G190), .A3(new_n551), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT83), .B1(new_n568), .B2(new_n571), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n568), .A2(KEYINPUT83), .A3(new_n571), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n554), .A2(G200), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n507), .A2(G68), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  INV_X1    g0383(.A(G97), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n350), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n206), .B1(new_n284), .B2(new_n583), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n404), .A2(new_n584), .A3(new_n359), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n247), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n520), .A2(G87), .A3(new_n521), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n351), .A2(new_n258), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G274), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n456), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n277), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT88), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(new_n277), .ZN(new_n599));
  INV_X1    g0399(.A(G250), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n205), .B2(G45), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n277), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT89), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n277), .A2(new_n604), .A3(new_n601), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n597), .A2(new_n599), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n280), .A2(G244), .A3(G1698), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n280), .A2(G238), .A3(new_n402), .ZN(new_n608));
  INV_X1    g0408(.A(new_n499), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n335), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n611), .A3(G190), .ZN(new_n612));
  INV_X1    g0412(.A(new_n599), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n598), .B1(new_n595), .B2(new_n277), .ZN(new_n614));
  INV_X1    g0414(.A(new_n605), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n604), .B1(new_n277), .B2(new_n601), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n613), .A2(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n499), .B1(new_n327), .B2(G238), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n277), .B1(new_n618), .B2(new_n607), .ZN(new_n619));
  OAI21_X1  g0419(.A(G200), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n593), .A2(new_n612), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n351), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n520), .A2(new_n623), .A3(new_n521), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n590), .A2(new_n624), .A3(new_n592), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G169), .B1(new_n617), .B2(new_n619), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n606), .A2(new_n611), .A3(G179), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT90), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n622), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n574), .A2(new_n581), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(G20), .B1(new_n252), .B2(G97), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n541), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G116), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G20), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(KEYINPUT20), .A3(new_n247), .A4(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n540), .B(KEYINPUT84), .ZN(new_n641));
  INV_X1    g0441(.A(new_n635), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n247), .A2(new_n638), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  MUX2_X1   g0446(.A(new_n257), .B(new_n519), .S(G116), .Z(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n280), .A2(G257), .A3(new_n402), .ZN(new_n649));
  INV_X1    g0449(.A(G303), .ZN(new_n650));
  INV_X1    g0450(.A(G264), .ZN(new_n651));
  OAI221_X1 g0451(.A(new_n649), .B1(new_n650), .B2(new_n280), .C1(new_n332), .C2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n301), .B1(new_n652), .B2(new_n335), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(G270), .B(new_n277), .C1(new_n474), .C2(new_n475), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n472), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n364), .B1(new_n646), .B2(new_n647), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n335), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n472), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT21), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT21), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n658), .A2(new_n663), .A3(new_n660), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n657), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n660), .A2(new_n305), .ZN(new_n667));
  INV_X1    g0467(.A(new_n648), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n660), .A2(G200), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n666), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n664), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n663), .B1(new_n658), .B2(new_n660), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n656), .B2(new_n654), .ZN(new_n674));
  INV_X1    g0474(.A(new_n670), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT91), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n634), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n453), .A2(new_n535), .A3(new_n677), .ZN(G372));
  NAND2_X1  g0478(.A1(new_n575), .A2(new_n551), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n555), .B1(new_n679), .B2(new_n364), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(new_n633), .A3(KEYINPUT26), .A4(new_n573), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n629), .A2(new_n625), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT83), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n566), .A2(new_n567), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n247), .ZN(new_n685));
  INV_X1    g0485(.A(new_n571), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n621), .B(new_n682), .C1(new_n687), .C2(new_n578), .ZN(new_n688));
  AOI21_X1  g0488(.A(G169), .B1(new_n575), .B2(new_n551), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(new_n555), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n681), .B1(new_n690), .B2(KEYINPUT26), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n492), .A2(new_n525), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n665), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n682), .A2(new_n621), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n528), .B2(new_n531), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n693), .A2(new_n574), .A3(new_n695), .A4(new_n581), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n691), .A2(new_n696), .A3(new_n682), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n453), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n346), .ZN(new_n699));
  INV_X1    g0499(.A(new_n311), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n366), .ZN(new_n701));
  INV_X1    g0501(.A(new_n304), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n447), .A2(KEYINPUT17), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT77), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n447), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT78), .B1(new_n447), .B2(KEYINPUT17), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n373), .B1(new_n441), .B2(new_n442), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n417), .A3(new_n444), .A4(new_n446), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n416), .B1(new_n703), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT99), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n712), .A2(new_n713), .B1(new_n340), .B2(new_n342), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n699), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n698), .A2(new_n716), .ZN(G369));
  NAND2_X1  g0517(.A1(new_n676), .A2(new_n671), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n265), .A2(new_n206), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT27), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT27), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G213), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G343), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n718), .B1(new_n668), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n674), .A2(new_n648), .A3(new_n724), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT100), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(G330), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n526), .A2(new_n725), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n525), .A2(new_n724), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n535), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n665), .A2(new_n724), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n535), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n492), .A2(new_n525), .A3(new_n725), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT101), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(KEYINPUT101), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n737), .A2(new_n745), .ZN(G399));
  INV_X1    g0546(.A(new_n209), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n289), .A2(new_n290), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n205), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n587), .A2(G116), .ZN(new_n753));
  INV_X1    g0553(.A(new_n750), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n752), .A2(new_n753), .B1(new_n215), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  INV_X1    g0556(.A(G330), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n677), .B(new_n725), .C1(new_n533), .C2(new_n534), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n617), .A2(new_n619), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G179), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n490), .A2(new_n760), .A3(new_n660), .A4(new_n554), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n653), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n656), .A3(new_n484), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n575), .A3(new_n551), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT30), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n763), .A2(KEYINPUT30), .A3(new_n575), .A4(new_n551), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n725), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT31), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n757), .B1(new_n758), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT26), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n680), .A2(new_n633), .A3(new_n772), .A4(new_n573), .ZN(new_n773));
  INV_X1    g0573(.A(new_n682), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n579), .A2(new_n577), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n682), .A2(new_n621), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n680), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(new_n777), .B2(KEYINPUT26), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n526), .A2(new_n665), .ZN(new_n779));
  AND3_X1   g0579(.A1(new_n579), .A2(new_n577), .A3(new_n580), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n576), .A2(new_n780), .B1(new_n680), .B2(new_n573), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n695), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n773), .B(new_n778), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(KEYINPUT102), .A3(new_n725), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(KEYINPUT102), .B1(new_n783), .B2(new_n725), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT29), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n697), .A2(new_n725), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT29), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n771), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n756), .B1(new_n791), .B2(G1), .ZN(G364));
  INV_X1    g0592(.A(new_n732), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n206), .A2(G13), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT103), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n751), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n729), .A2(new_n731), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G330), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G13), .A2(G33), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(G20), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n206), .A2(new_n301), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(G190), .A3(new_n309), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n280), .B1(new_n811), .B2(new_n349), .C1(new_n376), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n809), .A2(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n305), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G50), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n206), .A2(G179), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n818), .A2(G190), .A3(G200), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n816), .A2(new_n817), .B1(new_n819), .B2(new_n404), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n818), .A2(new_n305), .A3(G200), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n359), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n206), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n584), .ZN(new_n825));
  OR4_X1    g0625(.A1(new_n813), .A2(new_n820), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n818), .A2(new_n810), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT104), .B(G159), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT32), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n814), .A2(G190), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n262), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n819), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n815), .A2(G326), .B1(new_n834), .B2(G303), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n836), .B2(new_n821), .C1(new_n481), .C2(new_n824), .ZN(new_n837));
  INV_X1    g0637(.A(new_n812), .ZN(new_n838));
  INV_X1    g0638(.A(new_n827), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n838), .A2(G322), .B1(new_n839), .B2(G329), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT33), .B(G317), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(KEYINPUT105), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n831), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n811), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n280), .B1(new_n845), .B2(G311), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n840), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n826), .A2(new_n833), .B1(new_n837), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n213), .B1(G20), .B2(new_n364), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n806), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n747), .A2(new_n280), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(G45), .B2(new_n215), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n241), .B2(G45), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n747), .A2(new_n330), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(G355), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(G116), .B2(new_n209), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n851), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n850), .A2(new_n798), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n800), .A2(new_n803), .B1(new_n808), .B2(new_n859), .ZN(G396));
  INV_X1    g0660(.A(new_n828), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n838), .A2(G143), .B1(new_n845), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(new_n832), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G137), .B2(new_n815), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(KEYINPUT34), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(KEYINPUT34), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n280), .B1(new_n827), .B2(new_n868), .C1(new_n262), .C2(new_n821), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n824), .A2(new_n376), .B1(new_n819), .B2(new_n817), .ZN(new_n870));
  NOR4_X1   g0670(.A1(new_n866), .A2(new_n867), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n815), .A2(G303), .B1(new_n845), .B2(G116), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n836), .B2(new_n832), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT106), .Z(new_n874));
  AOI21_X1  g0674(.A(new_n825), .B1(G294), .B2(new_n838), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT107), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n821), .A2(new_n404), .ZN(new_n877));
  INV_X1    g0677(.A(G311), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n330), .B1(new_n827), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n877), .B(new_n879), .C1(G107), .C2(new_n834), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n874), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n849), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n849), .A2(new_n804), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n797), .B1(new_n349), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n366), .A2(new_n724), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n357), .A2(new_n724), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n369), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n366), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n882), .B(new_n884), .C1(new_n888), .C2(new_n805), .ZN(new_n889));
  INV_X1    g0689(.A(new_n771), .ZN(new_n890));
  INV_X1    g0690(.A(new_n888), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n788), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n366), .A2(new_n369), .A3(new_n725), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n697), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n798), .B1(new_n890), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n890), .A2(new_n896), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(G384));
  NOR2_X1   g0700(.A1(new_n563), .A2(new_n565), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n214), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT36), .Z(new_n906));
  OAI211_X1 g0706(.A(new_n216), .B(G77), .C1(new_n376), .C2(new_n218), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n817), .A2(G68), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n205), .B(G13), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n722), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n416), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT110), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n304), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n275), .B(KEYINPUT110), .C1(new_n302), .C2(new_n303), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n275), .A2(new_n724), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n915), .A2(new_n311), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n303), .ZN(new_n919));
  INV_X1    g0719(.A(new_n302), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n311), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n275), .A3(new_n724), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT109), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n885), .B(KEYINPUT108), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n895), .B2(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT109), .B(new_n925), .C1(new_n697), .C2(new_n894), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT16), .B1(new_n378), .B2(new_n390), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n374), .B1(new_n440), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n911), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n451), .B2(new_n416), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n398), .A2(new_n911), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT37), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n411), .A2(new_n935), .A3(new_n936), .A4(new_n447), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n931), .B1(new_n410), .B2(new_n911), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n447), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT37), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n933), .A2(new_n934), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n932), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n711), .B2(new_n415), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n913), .B1(new_n929), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT111), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n529), .A2(new_n530), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n776), .B1(new_n950), .B2(new_n525), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n665), .B2(new_n692), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n774), .B1(new_n952), .B2(new_n781), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n893), .B1(new_n953), .B2(new_n691), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT109), .B1(new_n954), .B2(new_n925), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n895), .A2(new_n924), .A3(new_n926), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n934), .B1(new_n933), .B2(new_n942), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n945), .A2(KEYINPUT38), .A3(new_n941), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n960), .A3(new_n923), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT111), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n913), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n949), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n915), .A2(new_n916), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n725), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT39), .B1(new_n943), .B2(new_n946), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT112), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n935), .B1(new_n451), .B2(new_n416), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n935), .A2(new_n411), .A3(new_n447), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(new_n936), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n934), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT39), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(new_n974), .A3(new_n959), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n969), .B1(new_n968), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n964), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n787), .A2(new_n453), .A3(new_n790), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n716), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT40), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n923), .A2(new_n888), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n758), .B2(new_n770), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n943), .B2(new_n946), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n973), .B2(new_n959), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n984), .A2(new_n987), .B1(new_n988), .B2(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n758), .A2(new_n770), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n453), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(G330), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n989), .B1(new_n453), .B2(new_n990), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n983), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n205), .B2(new_n795), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n983), .A2(new_n994), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n910), .B1(new_n996), .B2(new_n997), .ZN(G367));
  NOR2_X1   g0798(.A1(new_n593), .A2(new_n725), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n774), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n694), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n775), .A2(new_n724), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n680), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n781), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n574), .B1(new_n1007), .B2(new_n526), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n725), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n535), .A2(new_n738), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(KEYINPUT42), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1002), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n737), .A2(new_n1007), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n750), .B(KEYINPUT41), .Z(new_n1024));
  NAND2_X1  g0824(.A1(new_n745), .A2(new_n1006), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n745), .A2(new_n1006), .A3(new_n1026), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n743), .A2(new_n744), .A3(new_n1007), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT44), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n736), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT44), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1031), .B(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1035), .A2(new_n737), .A3(new_n1029), .A4(new_n1028), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n735), .B1(new_n665), .B2(new_n724), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n739), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(new_n793), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1033), .A2(new_n1036), .A3(new_n791), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1024), .B1(new_n1040), .B2(new_n791), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n796), .A2(G1), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1022), .B(new_n1023), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n852), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n851), .B1(new_n209), .B2(new_n351), .C1(new_n1044), .C2(new_n236), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT115), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n797), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n812), .A2(new_n863), .B1(new_n811), .B2(new_n817), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n330), .B(new_n1049), .C1(G137), .C2(new_n839), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n834), .A2(G58), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n821), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n831), .A2(new_n861), .B1(new_n1052), .B2(G77), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n824), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G68), .A2(new_n1054), .B1(new_n815), .B2(G143), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n824), .A2(new_n359), .B1(new_n811), .B2(new_n836), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT116), .Z(new_n1058));
  INV_X1    g0858(.A(G317), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n330), .B1(new_n827), .B2(new_n1059), .C1(new_n812), .C2(new_n650), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n831), .A2(G294), .B1(new_n1052), .B2(G97), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n878), .B2(new_n816), .ZN(new_n1062));
  OR3_X1    g0862(.A1(new_n1058), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT117), .B1(new_n819), .B2(new_n637), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT46), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1056), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT47), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1048), .B1(new_n1067), .B2(new_n849), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n807), .B2(new_n1001), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1043), .A2(new_n1069), .ZN(G387));
  OAI22_X1  g0870(.A1(new_n811), .A2(new_n262), .B1(new_n827), .B2(new_n863), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n330), .B(new_n1071), .C1(G50), .C2(new_n838), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n834), .A2(G77), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n623), .A2(new_n1054), .B1(new_n831), .B2(new_n317), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n815), .A2(G159), .B1(new_n1052), .B2(G97), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n280), .B1(new_n839), .B2(G326), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n824), .A2(new_n836), .B1(new_n819), .B2(new_n481), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n838), .A2(G317), .B1(new_n845), .B2(G303), .ZN(new_n1079));
  INV_X1    g0879(.A(G322), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n816), .B2(new_n1080), .C1(new_n878), .C2(new_n832), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1077), .B1(new_n637), .B2(new_n821), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n849), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n855), .A2(new_n753), .B1(new_n359), .B2(new_n747), .ZN(new_n1090));
  AOI211_X1 g0890(.A(G45), .B(new_n753), .C1(G68), .C2(G77), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT118), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n347), .A2(new_n817), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT50), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1093), .A2(KEYINPUT50), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(G45), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n852), .B1(new_n233), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1090), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n797), .B1(new_n1099), .B2(new_n851), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1089), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n735), .B2(new_n806), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1039), .A2(new_n791), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n750), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1039), .A2(new_n791), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(G393));
  INV_X1    g0907(.A(new_n1030), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n737), .B1(new_n1108), .B2(new_n1035), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1030), .A2(new_n1032), .A3(new_n736), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1104), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n750), .A3(new_n1040), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n852), .A2(new_n244), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n851), .C1(new_n584), .C2(new_n209), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n330), .B1(new_n839), .B2(G143), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n404), .B2(new_n821), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n824), .A2(new_n349), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n218), .B2(new_n819), .C1(new_n817), .C2(new_n832), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1116), .B(new_n1119), .C1(new_n347), .C2(new_n845), .ZN(new_n1120));
  INV_X1    g0920(.A(G159), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n816), .A2(new_n863), .B1(new_n1121), .B2(new_n812), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n816), .A2(new_n1059), .B1(new_n878), .B2(new_n812), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT52), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n832), .A2(new_n650), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n330), .B1(new_n827), .B2(new_n1080), .C1(new_n481), .C2(new_n811), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n824), .A2(new_n637), .B1(new_n819), .B2(new_n836), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n822), .A4(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1120), .A2(new_n1123), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n849), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n798), .B(new_n1114), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT119), .Z(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1007), .B2(new_n806), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n1042), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1112), .A2(new_n1136), .ZN(G390));
  AND3_X1   g0937(.A1(new_n973), .A2(new_n974), .A3(new_n959), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n974), .B1(new_n958), .B2(new_n959), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT112), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n929), .A2(new_n966), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n976), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n967), .B1(new_n973), .B2(new_n959), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n783), .A2(new_n725), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT102), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n885), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n784), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n887), .A2(new_n366), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n923), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1143), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n771), .A2(new_n888), .A3(new_n923), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1142), .A2(new_n1154), .A3(new_n1152), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n453), .A2(new_n771), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n981), .A2(new_n716), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n923), .B1(new_n771), .B2(new_n888), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1150), .A2(new_n1163), .A3(new_n1154), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n957), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1161), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n754), .B1(new_n1158), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1165), .B2(new_n1164), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1156), .A2(new_n1157), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1156), .A2(new_n1042), .A3(new_n1157), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n883), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n798), .B1(new_n317), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n812), .A2(new_n868), .B1(new_n811), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n330), .B(new_n1176), .C1(G125), .C2(new_n839), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n819), .A2(new_n863), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n831), .A2(G137), .B1(new_n1052), .B2(G50), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n824), .A2(new_n1121), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G128), .B2(new_n815), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n815), .A2(G283), .B1(new_n845), .B2(G97), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n359), .B2(new_n832), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  OAI221_X1 g0986(.A(new_n330), .B1(new_n827), .B2(new_n481), .C1(new_n812), .C2(new_n637), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n262), .A2(new_n821), .B1(new_n819), .B2(new_n404), .ZN(new_n1188));
  OR3_X1    g0988(.A1(new_n1187), .A2(new_n1117), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1183), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1174), .B1(new_n1190), .B2(new_n849), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n977), .A2(new_n978), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1193), .B2(new_n805), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1172), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT121), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1172), .B2(new_n1194), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1171), .B1(new_n1196), .B2(new_n1198), .ZN(G378));
  AOI21_X1  g0999(.A(new_n1151), .B1(new_n955), .B2(new_n956), .ZN(new_n1200));
  AOI211_X1 g1000(.A(KEYINPUT111), .B(new_n912), .C1(new_n1200), .C2(new_n960), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n962), .B1(new_n961), .B2(new_n913), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n966), .B1(new_n1140), .B2(new_n976), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n343), .A2(new_n346), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n322), .A2(new_n911), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n989), .B2(G330), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n987), .A2(new_n984), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n988), .A2(new_n986), .ZN(new_n1212));
  AND4_X1   g1012(.A1(G330), .A2(new_n1211), .A3(new_n1212), .A4(new_n1209), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1203), .A2(new_n1204), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(G330), .A3(new_n1212), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1209), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n989), .A2(G330), .A3(new_n1209), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n964), .A2(new_n979), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT123), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n980), .B(KEYINPUT123), .C1(new_n1213), .C2(new_n1210), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1042), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n797), .B1(new_n817), .B2(new_n883), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n839), .C2(G124), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n821), .B2(new_n828), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n815), .A2(G125), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n832), .B2(new_n868), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n838), .A2(G128), .B1(new_n845), .B2(G137), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n819), .B2(new_n1175), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G150), .C2(new_n1054), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1226), .B1(new_n1232), .B2(KEYINPUT59), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(KEYINPUT59), .B2(new_n1232), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n816), .A2(new_n637), .B1(new_n821), .B2(new_n376), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G97), .B2(new_n831), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n280), .B(new_n749), .C1(G283), .C2(new_n839), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n838), .A2(G107), .B1(new_n845), .B2(new_n623), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1054), .A2(G68), .B1(new_n834), .B2(G77), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n817), .B1(G33), .B2(G41), .C1(new_n749), .C2(new_n280), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1244));
  AND4_X1   g1044(.A1(new_n1234), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1224), .B1(new_n1131), .B2(new_n1245), .C1(new_n1209), .C2(new_n805), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1223), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1142), .A2(new_n1154), .A3(new_n1152), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1154), .B1(new_n1142), .B2(new_n1152), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1160), .B1(new_n1253), .B2(new_n1166), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1249), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1170), .A2(new_n1161), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1249), .B1(new_n1214), .B2(new_n1219), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n754), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1248), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(G375));
  INV_X1    g1060(.A(new_n1024), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1160), .A2(new_n1165), .A3(new_n1164), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1167), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1151), .A2(new_n804), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n637), .A2(new_n832), .B1(new_n816), .B2(new_n481), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G97), .B2(new_n834), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1052), .A2(G77), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1054), .A2(new_n623), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n812), .A2(new_n836), .B1(new_n811), .B2(new_n359), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n280), .B(new_n1269), .C1(G303), .C2(new_n839), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n824), .A2(new_n817), .B1(new_n819), .B2(new_n1121), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G132), .B2(new_n815), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n330), .B1(new_n839), .B2(G128), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n838), .A2(G137), .B1(new_n845), .B2(G150), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1175), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n831), .A2(new_n1276), .B1(new_n1052), .B2(G58), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1131), .B1(new_n1271), .B2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n797), .B(new_n1279), .C1(new_n262), .C2(new_n883), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1166), .A2(new_n1042), .B1(new_n1264), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1263), .A2(new_n1281), .ZN(G381));
  INV_X1    g1082(.A(G396), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G387), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1195), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1259), .A4(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1259), .A2(new_n1287), .A3(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(G407), .A2(G213), .A3(new_n1291), .ZN(G409));
  NAND2_X1  g1092(.A1(G393), .A2(G396), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1284), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1112), .A2(new_n1136), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1112), .B2(new_n1136), .ZN(new_n1297));
  OAI21_X1  g1097(.A(G387), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1294), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1300), .A2(new_n1043), .A3(new_n1069), .A4(new_n1295), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT61), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1160), .A2(new_n1165), .A3(new_n1164), .A4(KEYINPUT60), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(KEYINPUT125), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1262), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n750), .B(new_n1167), .C1(new_n1306), .C2(KEYINPUT60), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1281), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(G384), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G384), .B(new_n1281), .C1(new_n1305), .C2(new_n1307), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1290), .A2(G2897), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1214), .A2(new_n1219), .A3(KEYINPUT124), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1042), .A3(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1256), .A2(new_n1261), .A3(new_n1222), .A4(new_n1221), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1247), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1259), .A2(G378), .B1(new_n1287), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1315), .B1(new_n1323), .B2(new_n1290), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1248), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(G378), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1322), .A2(new_n1287), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n1290), .B(new_n1325), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT62), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1303), .B(new_n1324), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1290), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1325), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1302), .B1(new_n1332), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT63), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1302), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1330), .A2(KEYINPUT63), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1340), .A2(new_n1303), .A3(new_n1341), .A4(new_n1324), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1338), .A2(new_n1342), .ZN(G405));
  NAND2_X1  g1143(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1298), .A2(new_n1301), .A3(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1287), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1328), .B(KEYINPUT126), .C1(new_n1259), .C2(new_n1347), .ZN(new_n1348));
  OR3_X1    g1148(.A1(new_n1259), .A2(KEYINPUT126), .A3(new_n1347), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1349), .A3(new_n1325), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1325), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1344), .B(new_n1346), .C1(new_n1351), .C2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1352), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1345), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1354), .A2(new_n1355), .A3(new_n1350), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1356), .ZN(G402));
endmodule


