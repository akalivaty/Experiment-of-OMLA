//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT76), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n188), .A2(KEYINPUT76), .A3(G125), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n187), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G237), .ZN(new_n199));
  INV_X1    g013(.A(G953), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G214), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(G237), .A2(G953), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n209), .A3(new_n205), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n194), .A2(new_n187), .A3(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n198), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT86), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n203), .A2(new_n220), .A3(new_n205), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT18), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n203), .A2(new_n220), .A3(new_n224), .A4(new_n205), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n189), .A2(new_n191), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n192), .A2(new_n193), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(new_n187), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n226), .A2(KEYINPUT87), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT87), .B1(new_n226), .B2(new_n231), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n214), .B(new_n219), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n231), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n231), .A3(KEYINPUT87), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n230), .A2(KEYINPUT19), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT19), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(G146), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT88), .B1(new_n243), .B2(new_n197), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n207), .A2(new_n210), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n192), .B2(new_n193), .ZN(new_n246));
  INV_X1    g060(.A(new_n242), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n187), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n198), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n239), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n234), .B1(new_n252), .B2(new_n217), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(KEYINPUT90), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n217), .B1(new_n239), .B2(new_n251), .ZN(new_n257));
  INV_X1    g071(.A(new_n234), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n254), .B(new_n255), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT20), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n256), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G475), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n211), .A2(new_n213), .ZN(new_n266));
  INV_X1    g080(.A(new_n212), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(new_n197), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n237), .A2(new_n238), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n234), .B1(new_n269), .B2(new_n217), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT91), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n264), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n278));
  INV_X1    g092(.A(G122), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G116), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G122), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G107), .ZN(new_n284));
  XNOR2_X1  g098(.A(G116), .B(G122), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n278), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(G128), .B(G143), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n202), .A2(G128), .ZN(new_n291));
  OAI21_X1  g105(.A(G134), .B1(new_n291), .B2(KEYINPUT13), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n289), .B(G134), .C1(KEYINPUT13), .C2(new_n291), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(G107), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n286), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT92), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(KEYINPUT14), .A3(G122), .ZN(new_n300));
  OAI211_X1 g114(.A(G107), .B(new_n300), .C1(new_n283), .C2(KEYINPUT14), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n290), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n289), .A2(G134), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n297), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G217), .A3(new_n200), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT94), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n312), .A3(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT93), .B1(new_n306), .B2(new_n309), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n316));
  INV_X1    g130(.A(new_n309), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n299), .A2(new_n316), .A3(new_n305), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n271), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n311), .A2(new_n313), .B1(new_n315), .B2(new_n318), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT95), .B1(new_n323), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(G478), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(KEYINPUT15), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n320), .B(new_n271), .C1(KEYINPUT15), .C2(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G234), .A2(G237), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G952), .A3(new_n200), .ZN(new_n331));
  XOR2_X1   g145(.A(new_n331), .B(KEYINPUT96), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT21), .B(G898), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n330), .A2(G902), .A3(G953), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n275), .A2(new_n277), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n286), .A3(G104), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n216), .A2(G107), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT80), .A4(new_n342), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n345), .A2(new_n346), .A3(G101), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n187), .A2(G143), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n202), .A2(G146), .ZN(new_n350));
  AND2_X1   g164(.A1(KEYINPUT0), .A2(G128), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G143), .B(G146), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G128), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n216), .A2(KEYINPUT3), .A3(G107), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n286), .A2(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  INV_X1    g175(.A(G101), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n339), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n339), .A2(new_n341), .A3(new_n362), .A4(new_n342), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n345), .A2(G101), .A3(new_n347), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(KEYINPUT4), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n202), .A2(G146), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n187), .A2(G143), .ZN(new_n371));
  OAI211_X1 g185(.A(G128), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G128), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n349), .B(new_n350), .C1(KEYINPUT1), .C2(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n286), .A2(G104), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n362), .B1(new_n376), .B2(new_n342), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n375), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n357), .A2(new_n368), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n366), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n372), .A2(new_n374), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n382), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT11), .B1(new_n302), .B2(G137), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT11), .ZN(new_n392));
  INV_X1    g206(.A(G137), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT65), .B1(new_n393), .B2(G134), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT65), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n302), .A3(G137), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n209), .A2(new_n395), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n396), .A2(new_n398), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n209), .B1(new_n400), .B2(new_n395), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n383), .A2(new_n390), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n384), .A2(new_n388), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n381), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n209), .A3(new_n395), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT12), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT12), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n411), .B(new_n402), .C1(new_n404), .C2(new_n381), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n403), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G140), .ZN(new_n414));
  INV_X1    g228(.A(G227), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G953), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n414), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n383), .A2(new_n390), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n409), .ZN(new_n420));
  INV_X1    g234(.A(new_n417), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n403), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT83), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n418), .A2(new_n425), .A3(new_n422), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(G469), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n383), .A2(new_n390), .A3(new_n402), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n402), .B1(new_n383), .B2(new_n390), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n417), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n403), .B(new_n421), .C1(new_n410), .C2(new_n412), .ZN(new_n431));
  AOI211_X1 g245(.A(G469), .B(G902), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n271), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G221), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n308), .B2(new_n271), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G214), .B1(G237), .B2(G902), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G210), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT82), .B1(new_n366), .B2(new_n378), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n385), .B(new_n377), .C1(new_n363), .C2(new_n365), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT68), .B1(new_n281), .B2(G119), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT68), .ZN(new_n450));
  INV_X1    g264(.A(G119), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n281), .A2(G119), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT2), .ZN(new_n457));
  INV_X1    g271(.A(G113), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n459), .A2(new_n460), .B1(new_n457), .B2(new_n458), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n449), .A2(new_n452), .A3(KEYINPUT5), .A4(new_n453), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n281), .A2(KEYINPUT5), .A3(G119), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n458), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n455), .A2(new_n461), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n447), .A2(new_n448), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n455), .B(new_n461), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n368), .A2(new_n468), .A3(new_n348), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n446), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n386), .A2(new_n465), .A3(new_n387), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n368), .A2(new_n468), .A3(new_n348), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n445), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n446), .C1(new_n467), .C2(new_n469), .ZN(new_n476));
  AOI21_X1  g290(.A(G125), .B1(new_n372), .B2(new_n374), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n477), .A2(new_n478), .B1(G125), .B2(new_n355), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT84), .B1(new_n375), .B2(G125), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G224), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n481), .B(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n474), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT7), .B1(new_n482), .B2(G953), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n486), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n445), .B(KEYINPUT8), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n366), .A2(new_n465), .A3(new_n378), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n465), .B1(new_n366), .B2(new_n378), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT85), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n487), .A3(KEYINPUT85), .A4(new_n489), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n473), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n271), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n444), .B1(new_n485), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n497), .A2(new_n473), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  INV_X1    g316(.A(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n490), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n474), .A2(new_n476), .A3(new_n484), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n443), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n442), .B1(new_n500), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n338), .A2(new_n440), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n356), .B1(new_n399), .B2(new_n401), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n461), .B(new_n454), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n302), .A2(G137), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n393), .A2(G134), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n375), .A2(new_n408), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n468), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT72), .B1(new_n523), .B2(KEYINPUT28), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n204), .A2(G210), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT27), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(G101), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT29), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n528), .A2(new_n529), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT64), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n355), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n352), .B(KEYINPUT64), .C1(new_n353), .C2(new_n354), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT66), .B1(new_n402), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT66), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n409), .A2(new_n542), .A3(new_n538), .A4(new_n539), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n543), .A3(new_n517), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n468), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n518), .A2(new_n525), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n526), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n533), .B(KEYINPUT70), .Z(new_n548));
  OAI21_X1  g362(.A(new_n536), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n512), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n468), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n533), .B1(new_n554), .B2(new_n518), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n271), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G472), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n513), .B(new_n552), .C1(new_n544), .C2(new_n550), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n518), .A2(new_n533), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n561), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(KEYINPUT69), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(KEYINPUT31), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n552), .B1(new_n544), .B2(new_n550), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n566), .B2(new_n468), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n567), .A2(new_n568), .B1(new_n547), .B2(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT32), .B(new_n573), .C1(new_n565), .C2(new_n569), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n557), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT74), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n557), .B(new_n577), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  XOR2_X1   g392(.A(G119), .B(G128), .Z(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT23), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n451), .B2(G128), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n373), .A2(KEYINPUT23), .A3(G119), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n584), .C1(G119), .C2(new_n373), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n581), .B1(new_n585), .B2(G110), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n581), .B(new_n588), .C1(G110), .C2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n197), .A2(new_n228), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n579), .A2(new_n580), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(G110), .B2(new_n585), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n267), .B2(new_n197), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(KEYINPUT78), .A3(new_n595), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT22), .B(G137), .ZN(new_n600));
  INV_X1    g414(.A(G234), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n437), .A2(new_n601), .A3(G953), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n600), .B(new_n602), .Z(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n597), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n271), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT25), .ZN(new_n609));
  OAI21_X1  g423(.A(G217), .B1(new_n601), .B2(G902), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT75), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n605), .B2(new_n606), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT25), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n611), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(G902), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n609), .A2(new_n614), .B1(new_n607), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n576), .A2(new_n578), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n578), .A4(new_n617), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n511), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(new_n362), .ZN(G3));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n275), .A2(new_n277), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n309), .A2(KEYINPUT98), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n306), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n306), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(KEYINPUT33), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n323), .B2(KEYINPUT33), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n271), .A2(G478), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n624), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n264), .A2(new_n276), .A3(new_n273), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n276), .B1(new_n264), .B2(new_n273), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n624), .B(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n570), .A2(new_n571), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n565), .B2(new_n569), .ZN(new_n642));
  INV_X1    g456(.A(G472), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT97), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  INV_X1    g461(.A(new_n617), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n440), .A2(new_n509), .A3(new_n648), .A4(new_n336), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n640), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI21_X1  g466(.A(new_n272), .B1(new_n263), .B2(new_n259), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n329), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n647), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  XOR2_X1   g471(.A(new_n596), .B(KEYINPUT100), .Z(new_n658));
  NOR2_X1   g472(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n596), .B(KEYINPUT100), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(KEYINPUT36), .B2(new_n604), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n662), .A3(new_n616), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n599), .A2(new_n604), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT78), .B1(new_n592), .B2(new_n595), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n606), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n613), .B(new_n271), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n615), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n612), .A2(new_n613), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n647), .A2(new_n510), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AND4_X1   g488(.A1(new_n508), .A2(new_n436), .A3(new_n439), .A4(new_n671), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n335), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n332), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n654), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n576), .A2(new_n675), .A3(new_n681), .A4(new_n578), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XOR2_X1   g497(.A(new_n678), .B(KEYINPUT39), .Z(new_n684));
  NAND3_X1  g498(.A1(new_n436), .A2(new_n439), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n523), .A2(new_n548), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n562), .A2(new_n564), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n271), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n572), .B2(new_n574), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n671), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n625), .A2(new_n441), .A3(new_n329), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n504), .A2(new_n473), .A3(new_n497), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n271), .A2(new_n506), .A3(new_n443), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n443), .B1(new_n505), .B2(new_n506), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT38), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n686), .A2(new_n692), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n202), .ZN(G45));
  AND3_X1   g515(.A1(new_n576), .A2(new_n675), .A3(new_n578), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n633), .B(new_n679), .C1(new_n635), .C2(new_n636), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n625), .A2(new_n705), .A3(new_n633), .A4(new_n679), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT102), .B(G146), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G48));
  NOR2_X1   g524(.A1(new_n509), .A2(new_n336), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n634), .B2(new_n638), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n430), .A2(new_n431), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n433), .B1(new_n713), .B2(new_n271), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n432), .A3(new_n438), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n576), .A2(new_n578), .A3(new_n617), .A4(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT41), .B(G113), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND2_X1  g533(.A1(new_n711), .A2(new_n654), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n281), .ZN(G18));
  INV_X1    g536(.A(new_n338), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n508), .A2(new_n715), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n693), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n576), .A2(new_n723), .A3(new_n725), .A4(new_n578), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR2_X1   g541(.A1(new_n635), .A2(new_n636), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n508), .A2(new_n329), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n548), .B1(new_n528), .B2(new_n529), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n567), .A2(new_n568), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n565), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n571), .B(KEYINPUT103), .Z(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n648), .A3(new_n644), .ZN(new_n736));
  INV_X1    g550(.A(new_n715), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n336), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n730), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  INV_X1    g554(.A(new_n724), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n735), .A2(new_n693), .A3(new_n644), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n704), .A2(new_n706), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT104), .B(G125), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n743), .B(new_n744), .ZN(G27));
  XOR2_X1   g559(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n746));
  NOR2_X1   g560(.A1(new_n428), .A2(new_n417), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n747), .A2(new_n420), .B1(new_n413), .B2(new_n417), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n434), .B1(new_n748), .B2(G469), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n713), .A2(new_n433), .A3(new_n271), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n438), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n698), .A3(KEYINPUT105), .A4(new_n441), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n500), .A2(new_n441), .A3(new_n507), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n418), .A2(G469), .A3(new_n422), .ZN(new_n755));
  INV_X1    g569(.A(new_n434), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n439), .B1(new_n757), .B2(new_n432), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n753), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n752), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n576), .A2(new_n760), .A3(new_n578), .A4(new_n617), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n704), .A2(new_n706), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n746), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n575), .A2(KEYINPUT42), .A3(new_n617), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n707), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NOR2_X1   g581(.A1(new_n761), .A2(new_n680), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n302), .ZN(G36));
  AOI21_X1  g583(.A(KEYINPUT45), .B1(new_n424), .B2(new_n426), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n433), .B(new_n770), .C1(KEYINPUT45), .C2(new_n748), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n771), .A2(new_n772), .A3(new_n434), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n771), .B2(new_n434), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n750), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n439), .A3(new_n684), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n647), .A2(new_n693), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n728), .A2(new_n633), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n728), .A2(new_n781), .A3(new_n633), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT44), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n754), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n784), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n777), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND2_X1  g603(.A1(new_n775), .A2(new_n439), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT47), .Z(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n648), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n792), .B(new_n762), .C1(new_n576), .C2(new_n578), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  OR4_X1    g609(.A1(new_n442), .A2(new_n779), .A3(new_n438), .A4(new_n648), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT107), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT107), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n714), .A2(new_n432), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT49), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n691), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(new_n699), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n780), .A2(new_n333), .A3(new_n736), .A4(new_n782), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n699), .A2(new_n442), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n803), .A2(new_n737), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT50), .B1(new_n805), .B2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  OR4_X1    g621(.A1(KEYINPUT112), .A2(new_n803), .A3(new_n737), .A4(new_n804), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n780), .A2(new_n333), .A3(new_n782), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n715), .A3(new_n786), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n692), .A2(new_n333), .A3(new_n617), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n737), .A3(new_n754), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n625), .A2(new_n633), .ZN(new_n814));
  AOI22_X1  g628(.A1(new_n811), .A2(new_n742), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT113), .B1(new_n805), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n808), .B2(new_n806), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n803), .A2(new_n754), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n799), .A2(new_n439), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n821), .B1(new_n791), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n811), .A2(new_n575), .A3(new_n617), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n813), .A2(new_n640), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n200), .A2(G952), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT115), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n810), .A2(new_n715), .A3(new_n736), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n827), .B(new_n829), .C1(new_n509), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n826), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT109), .B1(new_n671), .B2(new_n678), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n609), .A2(new_n614), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n663), .A4(new_n679), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n841), .A2(new_n691), .A3(new_n751), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n702), .A2(new_n707), .B1(new_n730), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n743), .A2(new_n682), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT52), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n730), .A2(new_n691), .A3(new_n751), .A4(new_n841), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n576), .A2(new_n675), .A3(new_n578), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n762), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n743), .A2(new_n682), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n704), .A2(new_n706), .A3(new_n760), .A4(new_n742), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT108), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n329), .A2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n678), .B(new_n272), .C1(new_n263), .C2(new_n259), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT108), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n671), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n440), .A2(new_n858), .A3(new_n754), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n576), .A3(new_n578), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n853), .B(new_n860), .C1(new_n761), .C2(new_n680), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n625), .A2(new_n633), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n855), .A2(new_n857), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n625), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n647), .A2(new_n864), .A3(new_n649), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n672), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n622), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n726), .A2(new_n739), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n717), .A2(new_n721), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n852), .A2(new_n867), .A3(new_n766), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT110), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT53), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n622), .A2(new_n866), .ZN(new_n875));
  INV_X1    g689(.A(new_n861), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n869), .A3(new_n766), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(new_n843), .B2(new_n844), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n849), .A2(new_n850), .A3(new_n846), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n874), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n869), .A2(new_n766), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT53), .A3(new_n852), .A4(new_n867), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT110), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n873), .A2(new_n884), .A3(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT111), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n622), .A2(new_n861), .A3(new_n866), .A4(KEYINPUT111), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n869), .A2(KEYINPUT53), .A3(new_n766), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n889), .A2(new_n891), .B1(new_n870), .B2(new_n874), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n823), .B1(new_n820), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n816), .A2(new_n819), .A3(KEYINPUT114), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n836), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n802), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n200), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n892), .A2(new_n271), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT56), .B1(new_n906), .B2(G210), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n474), .A2(new_n476), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT117), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n484), .B(KEYINPUT55), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n907), .B2(new_n911), .ZN(G51));
  XNOR2_X1  g727(.A(new_n434), .B(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n620), .A2(new_n621), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n510), .ZN(new_n916));
  INV_X1    g730(.A(new_n866), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n876), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT111), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n717), .A2(new_n868), .ZN(new_n920));
  INV_X1    g734(.A(new_n721), .ZN(new_n921));
  AND4_X1   g735(.A1(KEYINPUT53), .A2(new_n920), .A3(new_n766), .A4(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n875), .A2(new_n886), .A3(new_n876), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(new_n922), .A3(new_n852), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n881), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n893), .B1(new_n924), .B2(new_n881), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n914), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n894), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(KEYINPUT118), .A3(new_n914), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n933), .A3(new_n713), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n906), .A2(new_n771), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n904), .B1(new_n934), .B2(new_n935), .ZN(G54));
  NAND4_X1  g750(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(new_n253), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT119), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT119), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  INV_X1    g754(.A(new_n253), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n904), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(G60));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  NOR2_X1   g759(.A1(new_n631), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n926), .B2(new_n927), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT120), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n932), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n631), .B1(new_n895), .B2(new_n945), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n905), .ZN(G63));
  AND2_X1   g767(.A1(new_n660), .A2(new_n662), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n925), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n925), .A2(KEYINPUT122), .A3(new_n954), .A4(new_n957), .ZN(new_n961));
  INV_X1    g775(.A(new_n607), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n892), .B2(new_n956), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n905), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT121), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(KEYINPUT61), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT61), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G66));
  INV_X1    g782(.A(new_n334), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n200), .B1(new_n969), .B2(G224), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n875), .A2(new_n869), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(new_n200), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n909), .B1(G898), .B2(new_n200), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT123), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n972), .B(new_n974), .ZN(G69));
  OAI21_X1  g789(.A(G953), .B1(new_n415), .B2(new_n676), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n730), .A2(new_n575), .A3(new_n617), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI22_X1  g794(.A1(new_n776), .A2(new_n980), .B1(new_n680), .B2(new_n761), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n791), .B2(new_n793), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n844), .A2(new_n708), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n788), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n200), .A3(new_n766), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n240), .A2(new_n242), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n566), .B(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n676), .B2(new_n200), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n978), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n983), .A2(new_n700), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT62), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n864), .B(KEYINPUT124), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n685), .A2(new_n754), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n994), .A2(new_n915), .A3(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n794), .A2(new_n993), .A3(new_n788), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n997), .A2(new_n200), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n991), .B1(new_n998), .B2(new_n988), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n976), .A2(new_n977), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT126), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n999), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  NAND3_X1  g819(.A1(new_n982), .A2(new_n766), .A3(new_n985), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(new_n971), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n554), .A2(new_n518), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1008), .A2(new_n533), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n904), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n873), .A2(new_n884), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n562), .A2(new_n564), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1011), .B(new_n1005), .C1(new_n1012), .C2(new_n555), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1005), .B1(new_n997), .B2(new_n971), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n533), .A3(new_n1008), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(G57));
endmodule


