//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  OR3_X1    g0029(.A1(KEYINPUT65), .A2(G58), .A3(G68), .ZN(new_n230));
  OAI21_X1  g0030(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(G50), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(G20), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g0036(.A1(new_n215), .A2(new_n228), .A3(new_n229), .A4(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G222), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(G223), .A3(G1698), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n235), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n235), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(G274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G41), .A2(G45), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT71), .B1(new_n282), .B2(G1), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n281), .A2(new_n274), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n279), .B1(G226), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n270), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n234), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G50), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n208), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(new_n296), .B2(new_n292), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT8), .B(G58), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n209), .A2(G33), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n209), .B2(new_n201), .ZN(new_n301));
  INV_X1    g0101(.A(G150), .ZN(new_n302));
  INV_X1    g0102(.A(G33), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n209), .A2(new_n303), .A3(KEYINPUT73), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G20), .B2(G33), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n294), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n286), .A2(G179), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT75), .B(G200), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n286), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n309), .B(KEYINPUT9), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n286), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT76), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n255), .A2(G232), .A3(new_n256), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n255), .A2(G238), .A3(G1698), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n322), .B(new_n323), .C1(new_n205), .C2(new_n255), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n268), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n284), .A2(G244), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n278), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n321), .B1(new_n327), .B2(G179), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n279), .B1(G244), .B2(new_n284), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n329), .A2(KEYINPUT76), .A3(new_n330), .A4(new_n325), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n299), .B(KEYINPUT74), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n304), .A2(new_n306), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT15), .B(G87), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n300), .B1(new_n209), .B2(new_n202), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n294), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n295), .A2(new_n340), .B1(new_n202), .B2(new_n292), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n339), .A2(new_n341), .B1(new_n327), .B2(new_n287), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n327), .A2(new_n313), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n329), .A2(G190), .A3(new_n325), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n339), .A3(new_n341), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G226), .A2(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G232), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(G1698), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n354), .B2(new_n255), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(new_n267), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n281), .A2(new_n274), .A3(G238), .A4(new_n283), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n278), .A4(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n358), .B(new_n278), .C1(new_n355), .C2(new_n267), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT13), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(new_n361), .A3(new_n316), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n300), .A2(new_n202), .B1(new_n209), .B2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n294), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT78), .B(new_n294), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT11), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT12), .ZN(new_n377));
  INV_X1    g0177(.A(G68), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n292), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT12), .B1(new_n291), .B2(G68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n378), .B1(new_n208), .B2(G20), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n295), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n374), .A2(new_n376), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT79), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n384), .B1(new_n373), .B2(KEYINPUT11), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT79), .B1(new_n389), .B2(new_n376), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n366), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(KEYINPUT79), .A3(new_n376), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT80), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n366), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n362), .A2(G169), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n359), .A2(new_n361), .A3(G179), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n362), .A2(new_n403), .A3(G169), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n320), .A2(new_n349), .A3(new_n398), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n255), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n378), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(G58), .B(G68), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n334), .A2(G159), .B1(new_n413), .B2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n261), .B2(new_n209), .ZN(new_n417));
  NOR4_X1   g0217(.A1(new_n259), .A2(new_n260), .A3(new_n409), .A4(G20), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT16), .A3(new_n414), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n420), .A3(new_n294), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n299), .B1(new_n208), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n295), .A2(new_n422), .B1(new_n292), .B2(new_n299), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n281), .A2(new_n274), .A3(new_n283), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n278), .B1(new_n424), .B2(new_n353), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT82), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT82), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n255), .A2(new_n429), .A3(G226), .A4(G1698), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n255), .A2(G223), .A3(new_n256), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n428), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n268), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n426), .A2(new_n434), .A3(new_n316), .ZN(new_n435));
  AOI21_X1  g0235(.A(G200), .B1(new_n426), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n421), .B(new_n423), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n421), .A2(new_n423), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n421), .A2(new_n442), .A3(new_n423), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n426), .A2(new_n434), .A3(G179), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n425), .B1(new_n268), .B2(new_n433), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n287), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n440), .A2(new_n441), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n440), .A2(new_n443), .A3(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT18), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n438), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n407), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n294), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n291), .C1(G1), .C2(new_n303), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G116), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n292), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(G20), .B1(G33), .B2(G283), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G33), .B2(new_n204), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n294), .C1(new_n209), .C2(G116), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n455), .B(new_n457), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G257), .A2(G1698), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n256), .A2(G264), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n255), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(new_n268), .C1(G303), .C2(new_n255), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n208), .A2(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n274), .A3(G274), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n276), .A2(G1), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n274), .A2(new_n478), .A3(G270), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n469), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n465), .A2(KEYINPUT21), .A3(G169), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n457), .B1(new_n453), .B2(new_n456), .ZN(new_n483));
  OR2_X1    g0283(.A1(new_n460), .A2(new_n461), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n462), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n480), .A2(G169), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n480), .A2(new_n330), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n465), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n480), .A2(G200), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n485), .B(new_n491), .C1(new_n316), .C2(new_n480), .ZN(new_n492));
  OAI211_X1 g0292(.A(G244), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G250), .A2(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT4), .A2(G244), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(G1698), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n255), .A2(new_n498), .B1(G33), .B2(G283), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n267), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n274), .A2(new_n478), .A3(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n474), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT84), .B1(new_n500), .B2(new_n502), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(G200), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n292), .A2(new_n204), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n453), .B2(new_n204), .ZN(new_n509));
  OAI21_X1  g0309(.A(G107), .B1(new_n417), .B2(new_n418), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n334), .A2(G77), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n206), .A3(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n204), .A2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n510), .B(new_n511), .C1(new_n516), .C2(new_n209), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n509), .B1(new_n517), .B2(new_n294), .ZN(new_n518));
  INV_X1    g0318(.A(new_n503), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n507), .B(new_n518), .C1(new_n316), .C2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n518), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n500), .A2(new_n502), .A3(G179), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n503), .A2(G169), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AND4_X1   g0326(.A1(new_n490), .A2(new_n492), .A3(new_n520), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n274), .A2(new_n478), .A3(G264), .ZN(new_n528));
  INV_X1    g0328(.A(G294), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n303), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G250), .A2(G1698), .ZN(new_n531));
  INV_X1    g0331(.A(G257), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n532), .B2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n530), .B1(new_n533), .B2(new_n255), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n474), .B(new_n528), .C1(new_n534), .C2(new_n267), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G169), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT90), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT91), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n535), .B2(new_n330), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n274), .A2(new_n478), .A3(G264), .ZN(new_n540));
  OR2_X1    g0340(.A1(G250), .A2(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(G1698), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n259), .C2(new_n260), .ZN(new_n543));
  INV_X1    g0343(.A(new_n530), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n267), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT91), .A3(G179), .A4(new_n474), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT90), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n535), .A2(new_n548), .A3(G169), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n537), .A2(new_n539), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n209), .A2(G107), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n290), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT89), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(KEYINPUT25), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n556), .B1(new_n554), .B2(new_n552), .C1(new_n453), .C2(new_n205), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT88), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT88), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n562));
  OR3_X1    g0362(.A1(new_n209), .A2(KEYINPUT23), .A3(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n209), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT22), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n255), .A2(new_n568), .A3(new_n209), .A4(G87), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n294), .B1(new_n570), .B2(KEYINPUT24), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT24), .ZN(new_n572));
  AOI211_X1 g0372(.A(new_n572), .B(new_n565), .C1(new_n567), .C2(new_n569), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n558), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n550), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n535), .A2(new_n363), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G190), .B2(new_n535), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(new_n558), .C1(new_n573), .C2(new_n571), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n255), .A2(G244), .A3(G1698), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n255), .A2(G238), .A3(new_n256), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n303), .C2(new_n456), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n268), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT85), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n470), .A2(new_n584), .A3(G250), .ZN(new_n585));
  AOI21_X1  g0385(.A(G274), .B1(KEYINPUT85), .B2(G250), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n470), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n274), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n583), .A2(G190), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT87), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n582), .A2(new_n268), .B1(new_n274), .B2(new_n587), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT19), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n209), .B1(new_n350), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(G87), .B2(new_n206), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n209), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n300), .B2(new_n204), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n294), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n336), .A2(new_n291), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT86), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n606), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n454), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n583), .A2(new_n588), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n313), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n594), .A2(new_n608), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n601), .B2(new_n603), .ZN(new_n613));
  AOI211_X1 g0413(.A(KEYINPUT86), .B(new_n602), .C1(new_n600), .C2(new_n294), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n337), .B2(new_n453), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n591), .A2(new_n330), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n615), .B(new_n616), .C1(G169), .C2(new_n591), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(new_n451), .A2(new_n527), .A3(new_n579), .A4(new_n618), .ZN(G372));
  NAND2_X1  g0419(.A1(new_n318), .A2(new_n319), .ZN(new_n620));
  INV_X1    g0420(.A(new_n438), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n398), .A2(new_n332), .A3(new_n342), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n406), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n446), .A2(new_n439), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n624), .B(KEYINPUT18), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n620), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n312), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT92), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n610), .A2(new_n629), .A3(new_n287), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT92), .B1(new_n591), .B2(G169), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n615), .A2(new_n616), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n608), .A2(new_n589), .A3(new_n609), .A4(new_n611), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n520), .A2(new_n526), .A3(new_n578), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n490), .A2(new_n575), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n518), .A2(new_n524), .A3(new_n522), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n612), .A2(KEYINPUT26), .A3(new_n638), .A4(new_n617), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n451), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n628), .A2(new_n645), .ZN(G369));
  INV_X1    g0446(.A(KEYINPUT95), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n290), .A2(new_n209), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n574), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n575), .A2(new_n578), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT94), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT94), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n575), .A2(new_n657), .A3(new_n578), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n653), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n575), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n647), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  AOI211_X1 g0463(.A(KEYINPUT95), .B(new_n661), .C1(new_n656), .C2(new_n658), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT93), .B1(new_n490), .B2(new_n492), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n485), .A2(new_n660), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n490), .A2(KEYINPUT93), .A3(new_n492), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n490), .A2(new_n668), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n671), .A2(G330), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n490), .A2(new_n653), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n663), .B2(new_n664), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n550), .A2(new_n574), .A3(new_n660), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(G399));
  NAND3_X1  g0478(.A1(new_n212), .A2(KEYINPUT96), .A3(new_n275), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT96), .B1(new_n212), .B2(new_n275), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n232), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n618), .A2(new_n640), .A3(new_n638), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n637), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n688), .B1(new_n691), .B2(new_n660), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n488), .A2(new_n503), .A3(new_n546), .A4(new_n591), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT98), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n591), .A2(new_n503), .A3(new_n546), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT98), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT30), .A4(new_n488), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n480), .A2(new_n330), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n591), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n610), .A2(KEYINPUT97), .A3(new_n330), .A4(new_n480), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n503), .B1(new_n474), .B2(new_n546), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n695), .B2(new_n694), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n653), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n527), .A2(new_n579), .A3(new_n618), .A4(new_n660), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G330), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n653), .B1(new_n637), .B2(new_n643), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n688), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n693), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n687), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(new_n289), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n208), .B1(new_n721), .B2(G45), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n683), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n673), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(G330), .B1(new_n671), .B2(new_n672), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n671), .A2(new_n672), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n212), .A2(new_n255), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n733), .A2(new_n734), .B1(G116), .B2(new_n212), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n250), .A2(new_n276), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n212), .A2(new_n261), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n233), .B2(new_n276), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n234), .B1(G20), .B2(new_n287), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n724), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n209), .A2(new_n316), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n313), .A2(new_n330), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(G303), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n261), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT102), .Z(new_n748));
  NOR2_X1   g0548(.A1(new_n209), .A2(G190), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n313), .A2(new_n330), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT101), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G283), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G329), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n330), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n744), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n749), .A2(new_n760), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n316), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n768), .A2(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n209), .B1(new_n753), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n765), .B(new_n773), .C1(G294), .C2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n748), .A2(new_n752), .A3(new_n759), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n204), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n767), .B2(G68), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n296), .B2(new_n771), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT100), .B(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n757), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT32), .Z(new_n783));
  INV_X1    g0583(.A(new_n745), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n784), .A2(G87), .ZN(new_n785));
  INV_X1    g0585(.A(G58), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n255), .B1(new_n763), .B2(new_n202), .C1(new_n786), .C2(new_n761), .ZN(new_n787));
  OR4_X1    g0587(.A1(new_n780), .A2(new_n783), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n751), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n205), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n777), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n743), .B1(new_n791), .B2(new_n740), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n725), .A2(new_n727), .B1(new_n732), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  NAND3_X1  g0594(.A1(new_n332), .A2(new_n342), .A3(new_n653), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT103), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n332), .A2(KEYINPUT103), .A3(new_n342), .A4(new_n653), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n339), .A2(new_n341), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n343), .B(new_n346), .C1(new_n800), .C2(new_n660), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n716), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n641), .A2(new_n642), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n574), .B2(new_n550), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n520), .A2(new_n526), .A3(new_n578), .A4(new_n634), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n632), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n802), .B(new_n660), .C1(new_n804), .C2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OR3_X1    g0610(.A1(new_n715), .A2(new_n803), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n715), .B1(new_n803), .B2(new_n810), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n811), .A2(new_n723), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n740), .A2(new_n729), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n724), .B1(G77), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n771), .A2(new_n746), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n778), .B(new_n817), .C1(G283), .C2(new_n767), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n261), .B1(new_n763), .B2(new_n456), .C1(new_n529), .C2(new_n761), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G107), .B2(new_n784), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n751), .A2(G87), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n758), .A2(G311), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n761), .ZN(new_n824));
  INV_X1    g0624(.A(new_n763), .ZN(new_n825));
  INV_X1    g0625(.A(new_n781), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n824), .A2(G143), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n302), .B2(new_n768), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G137), .B2(new_n770), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n255), .B1(new_n774), .B2(new_n786), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n758), .B2(G132), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n751), .A2(G68), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n833), .C1(new_n296), .C2(new_n745), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n823), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n816), .B1(new_n835), .B2(new_n740), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n802), .B2(new_n730), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n813), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT104), .B1(new_n813), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G384));
  AND3_X1   g0641(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n842));
  INV_X1    g0642(.A(new_n397), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n396), .B1(new_n395), .B2(new_n366), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n395), .A2(new_n660), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT105), .B1(new_n842), .B2(new_n395), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT105), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n399), .A2(new_n405), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n846), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n398), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(new_n714), .A3(new_n802), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n421), .A2(new_n423), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n651), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n450), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n437), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n651), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n440), .A2(new_n443), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n861), .A2(new_n448), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n624), .A2(new_n437), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT106), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n624), .A2(new_n437), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n858), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n864), .B1(new_n870), .B2(KEYINPUT37), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n856), .B1(new_n859), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n861), .A2(new_n448), .A3(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n450), .A2(new_n858), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n872), .A2(KEYINPUT107), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT107), .B1(new_n872), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n855), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n863), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n621), .B2(new_n625), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT37), .B1(new_n883), .B2(new_n865), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n874), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n856), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n881), .B1(new_n888), .B2(new_n877), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n855), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n451), .A2(new_n714), .ZN(new_n893));
  OAI21_X1  g0693(.A(G330), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n872), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n848), .A2(new_n850), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n660), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT39), .B1(new_n888), .B2(new_n877), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n897), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n343), .A2(new_n653), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n809), .A2(new_n905), .B1(new_n847), .B2(new_n852), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n878), .B2(new_n879), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n625), .A2(new_n651), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n717), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n451), .B1(new_n910), .B2(new_n692), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n627), .A3(new_n626), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n909), .B(new_n912), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n895), .A2(new_n913), .B1(new_n208), .B2(new_n721), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n895), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n234), .A2(new_n209), .A3(new_n456), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT35), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n916), .B1(new_n516), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n917), .B2(new_n516), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n233), .B(G77), .C1(new_n786), .C2(new_n378), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n296), .A2(G68), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n208), .B(G13), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n915), .A2(new_n920), .A3(new_n923), .ZN(G367));
  NAND2_X1  g0724(.A1(new_n608), .A2(new_n609), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n633), .A2(new_n925), .A3(new_n653), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n653), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n632), .A3(new_n634), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n731), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n246), .A2(new_n212), .A3(new_n261), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n741), .C1(new_n212), .C2(new_n337), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT112), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n723), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  INV_X1    g0736(.A(new_n750), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n758), .A2(G137), .B1(new_n937), .B2(G77), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n786), .B2(new_n745), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n825), .A2(G50), .B1(new_n826), .B2(new_n767), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT113), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n774), .A2(new_n378), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n261), .B(new_n943), .C1(G150), .C2(new_n824), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n940), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n770), .A2(G143), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(G283), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n261), .B1(new_n763), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G303), .B2(new_n824), .ZN(new_n950));
  INV_X1    g0750(.A(G317), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n950), .B1(new_n204), .B2(new_n750), .C1(new_n951), .C2(new_n757), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n775), .A2(G107), .B1(G311), .B2(new_n770), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT46), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n745), .B2(new_n456), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n767), .A2(G294), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n953), .A2(new_n954), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n939), .A2(new_n947), .B1(new_n952), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT47), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n936), .B1(new_n960), .B2(new_n740), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n931), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT111), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n520), .B(new_n526), .C1(new_n518), .C2(new_n660), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n638), .A2(new_n653), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n676), .A2(new_n677), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n677), .A4(new_n966), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n676), .A2(new_n677), .ZN(new_n972));
  INV_X1    g0772(.A(new_n966), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT44), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n975), .B(new_n966), .C1(new_n676), .C2(new_n677), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n969), .A2(new_n971), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n674), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(new_n968), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n674), .C1(new_n974), .C2(new_n976), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n665), .B1(new_n490), .B2(new_n653), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n673), .A3(new_n676), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n673), .B1(new_n983), .B2(new_n676), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n985), .A2(new_n986), .A3(new_n718), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(new_n719), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n682), .B(KEYINPUT41), .Z(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT109), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n990), .B1(new_n988), .B2(new_n719), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n722), .B(KEYINPUT110), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n675), .B(new_n966), .C1(new_n663), .C2(new_n664), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n520), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n526), .B1(new_n1001), .B2(new_n575), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1000), .A2(KEYINPUT42), .B1(new_n660), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n998), .B(KEYINPUT108), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT42), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT43), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n930), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n978), .A2(new_n966), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1003), .A2(new_n1008), .A3(new_n930), .A4(new_n1006), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n963), .B1(new_n997), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n1019));
  AOI211_X1 g0819(.A(KEYINPUT109), .B(new_n990), .C1(new_n988), .C2(new_n719), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n963), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n962), .B1(new_n1018), .B2(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(KEYINPUT114), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n987), .B2(new_n683), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n986), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(new_n719), .A3(new_n984), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(KEYINPUT114), .A3(new_n682), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n718), .B1(new_n985), .B2(new_n986), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n261), .B1(new_n757), .B2(new_n772), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n824), .B1(new_n825), .B2(G303), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n771), .B2(new_n762), .C1(new_n764), .C2(new_n768), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT48), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n784), .A2(G294), .B1(G283), .B2(new_n775), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT49), .Z(new_n1039));
  AOI211_X1 g0839(.A(new_n1031), .B(new_n1039), .C1(G116), .C2(new_n937), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n775), .A2(new_n336), .ZN(new_n1041));
  INV_X1    g0841(.A(G159), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1041), .B1(new_n771), .B2(new_n1042), .C1(new_n299), .C2(new_n768), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n255), .B1(new_n761), .B2(new_n296), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G68), .B2(new_n825), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n784), .A2(G77), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n302), .C2(new_n757), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1043), .B(new_n1047), .C1(G97), .C2(new_n751), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n740), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n733), .A2(new_n684), .B1(G107), .B2(new_n212), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n333), .A2(new_n296), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT50), .Z(new_n1052));
  AOI21_X1  g0852(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n684), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n737), .B1(new_n243), .B2(G45), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1049), .B(new_n724), .C1(new_n742), .C2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n665), .B2(new_n731), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n985), .A2(new_n986), .A3(new_n996), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1030), .A2(new_n1060), .ZN(G393));
  NAND2_X1  g0861(.A1(new_n979), .A2(new_n982), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n996), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n973), .A2(new_n731), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n741), .B1(new_n204), .B2(new_n212), .C1(new_n253), .C2(new_n737), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n724), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n771), .A2(new_n302), .B1(new_n761), .B2(new_n1042), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT51), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n775), .A2(G77), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n255), .C1(new_n296), .C2(new_n768), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n758), .A2(G143), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n333), .A2(new_n825), .B1(new_n784), .B2(G68), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1073), .A2(new_n821), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n261), .B1(new_n757), .B2(new_n762), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1077), .B(new_n790), .C1(G283), .C2(new_n784), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT116), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n771), .A2(new_n951), .B1(new_n761), .B2(new_n764), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n767), .A2(G303), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n825), .A2(G294), .B1(new_n775), .B2(G116), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1066), .B1(new_n1086), .B2(new_n740), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1063), .B1(new_n1064), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1062), .A2(new_n1027), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n682), .A3(new_n988), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(G390));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n906), .B2(new_n900), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n904), .B1(new_n716), .B2(new_n802), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n847), .A2(new_n852), .ZN(new_n1095));
  OAI211_X1 g0895(.A(KEYINPUT118), .B(new_n899), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(new_n896), .C2(new_n901), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n899), .B(KEYINPUT117), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n888), .A2(new_n877), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n691), .A2(new_n660), .A3(new_n802), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n905), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1098), .B(new_n1099), .C1(new_n1101), .C2(new_n1095), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1097), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n714), .A2(G330), .A3(new_n802), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n1095), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1104), .A2(new_n1095), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1097), .A2(new_n1107), .A3(new_n1102), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n730), .B1(new_n897), .B2(new_n902), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n833), .B1(new_n529), .B2(new_n757), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT120), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1070), .B1(new_n771), .B2(new_n948), .C1(new_n205), .C2(new_n768), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n261), .B1(new_n763), .B2(new_n204), .C1(new_n456), .C2(new_n761), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1112), .A2(new_n785), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n261), .B1(new_n824), .B2(G132), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n763), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G50), .B2(new_n937), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n758), .A2(G125), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n767), .A2(G137), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n775), .A2(G159), .B1(G128), .B2(new_n770), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n745), .B2(new_n302), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n784), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n740), .B1(new_n1115), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n723), .B1(new_n299), .B2(new_n814), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1109), .A2(new_n996), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n451), .A2(G330), .A3(new_n714), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n628), .A2(new_n911), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1104), .A2(new_n1095), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT119), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1104), .A2(new_n1136), .A3(new_n1095), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1135), .A2(new_n1107), .A3(new_n1101), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1134), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1139), .A2(new_n1105), .B1(new_n810), .B2(new_n904), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1133), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n683), .B1(new_n1109), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1106), .A2(new_n1141), .A3(new_n1108), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1131), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(new_n1133), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT107), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n859), .A2(new_n871), .A3(new_n856), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT38), .B1(new_n875), .B2(new_n876), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT107), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n854), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n890), .C1(new_n1154), .C2(KEYINPUT40), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n309), .A2(new_n862), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n320), .B(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n909), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n882), .A2(G330), .A3(new_n890), .A4(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1161), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1148), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1148), .B(KEYINPUT57), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n682), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n909), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n996), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1159), .A2(new_n729), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n724), .B1(G50), .B2(new_n815), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n825), .A2(new_n336), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n255), .A2(G41), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n824), .A2(G107), .ZN(new_n1179));
  AND4_X1   g0979(.A1(new_n1046), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n771), .A2(new_n456), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n943), .B(new_n1181), .C1(G97), .C2(new_n767), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n758), .A2(G283), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n937), .A2(G58), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n296), .B1(G33), .B2(G41), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1185), .A2(new_n1186), .B1(new_n1178), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1186), .B2(new_n1185), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n824), .B1(new_n825), .B2(G137), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n745), .A2(new_n1117), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n767), .A2(G132), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n775), .A2(G150), .B1(G125), .B2(new_n770), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT59), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n303), .B(new_n275), .C1(new_n750), .C2(new_n781), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n758), .B2(G124), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1189), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1176), .B1(new_n1201), .B2(new_n740), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1174), .B1(new_n1175), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1170), .A2(new_n1203), .ZN(G375));
  AND3_X1   g1004(.A1(new_n1138), .A2(new_n1133), .A3(new_n1140), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1205), .A2(new_n1141), .A3(new_n990), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1095), .A2(new_n729), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT122), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n724), .B1(G68), .B2(new_n815), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1041), .B1(new_n771), .B2(new_n529), .C1(new_n456), .C2(new_n768), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n757), .A2(new_n746), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n745), .A2(new_n204), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n261), .B1(new_n763), .B2(new_n205), .C1(new_n948), .C2(new_n761), .ZN(new_n1213));
  OR4_X1    g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n789), .A2(new_n202), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n758), .A2(G128), .B1(G159), .B2(new_n784), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n255), .B1(new_n763), .B2(new_n302), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G137), .B2(new_n824), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1218), .A3(new_n1184), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n775), .A2(G50), .B1(G132), .B2(new_n770), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n768), .B2(new_n1117), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1214), .A2(new_n1215), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1209), .B1(new_n1222), .B2(new_n740), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1208), .A2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n996), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1206), .A2(new_n1226), .ZN(G381));
  NAND3_X1  g1027(.A1(new_n1030), .A2(new_n793), .A3(new_n1060), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(G384), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT123), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1230), .A2(G378), .A3(G390), .A4(G381), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n962), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT111), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1021), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1231), .A2(new_n1235), .A3(new_n1170), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n1145), .A2(new_n652), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G375), .C2(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(G343), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1138), .A2(new_n1133), .A3(new_n1140), .A4(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n682), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT60), .B1(new_n1225), .B2(new_n1133), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1205), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n840), .B1(new_n1246), .B2(new_n1226), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1226), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1205), .B1(new_n1142), .B2(KEYINPUT60), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G384), .B(new_n1248), .C1(new_n1249), .C2(new_n1243), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1241), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1241), .ZN(new_n1254));
  AOI211_X1 g1054(.A(KEYINPUT125), .B(new_n1254), .C1(new_n1247), .C2(new_n1250), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1253), .A2(new_n1255), .B1(new_n1252), .B2(new_n1251), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1170), .A2(G378), .A3(new_n1203), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT124), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1172), .A2(new_n1260), .A3(new_n1173), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1259), .A2(new_n1261), .A3(new_n995), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1175), .A2(new_n1202), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1166), .B2(new_n990), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1145), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1258), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1240), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT61), .B1(new_n1257), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1251), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1266), .A2(new_n1270), .A3(new_n1267), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1228), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n1090), .A3(new_n1088), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G390), .A2(new_n1228), .A3(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G387), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1276), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1279), .B1(new_n1235), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1240), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1270), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1269), .A2(new_n1273), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1280), .B1(G387), .B2(new_n1276), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1235), .A2(new_n1282), .A3(new_n1279), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1281), .A2(new_n1283), .A3(KEYINPUT127), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1285), .B2(new_n1256), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1271), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1285), .A2(KEYINPUT62), .A3(new_n1270), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1295), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1287), .B1(new_n1293), .B2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1145), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1258), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1270), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1251), .A3(new_n1258), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1305), .B(new_n1306), .ZN(G402));
endmodule


