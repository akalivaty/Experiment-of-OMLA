//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT65), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT66), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n474), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n460), .B2(G114), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  AOI211_X1 g071(.A(new_n496), .B(new_n489), .C1(new_n491), .C2(new_n493), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n474), .A2(KEYINPUT67), .A3(G126), .A4(G2105), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT70), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n475), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G138), .C1(new_n465), .C2(new_n466), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n501), .A2(new_n502), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n510), .B(new_n511), .C1(new_n495), .C2(new_n497), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n504), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT71), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(KEYINPUT5), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n524), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G88), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n529), .B1(new_n528), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n520), .B1(new_n536), .B2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n521), .A2(new_n523), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n516), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n526), .A2(G51), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n542), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n552), .B1(new_n543), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n515), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(G171));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT74), .B(G43), .Z(new_n559));
  OAI22_X1  g134(.A1(new_n558), .A2(new_n543), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n515), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G188));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  INV_X1    g146(.A(G78), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n533), .A2(new_n571), .B1(new_n572), .B2(new_n525), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI221_X1 g150(.A(KEYINPUT76), .B1(new_n572), .B2(new_n525), .C1(new_n533), .C2(new_n571), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(G651), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n534), .A2(G91), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n526), .B2(G53), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n526), .A2(new_n579), .A3(G53), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n577), .B(new_n578), .C1(new_n580), .C2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  NAND2_X1  g158(.A1(new_n526), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n542), .A2(G87), .A3(new_n516), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n533), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n526), .B2(G48), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n542), .A2(G86), .A3(new_n516), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n534), .A2(new_n594), .A3(G86), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(G305));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(new_n552), .B1(new_n543), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n515), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G171), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT78), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n542), .A2(G92), .A3(new_n516), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n526), .A2(G54), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n515), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(G868), .B2(new_n612), .ZN(G284));
  OAI21_X1  g188(.A(new_n606), .B1(G868), .B2(new_n612), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n604), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G168), .B2(new_n604), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(G168), .B2(new_n604), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n612), .B1(new_n618), .B2(G860), .ZN(G148));
  OR2_X1    g194(.A1(new_n560), .A2(new_n562), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n604), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n618), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n621), .B1(new_n623), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g200(.A1(new_n465), .A2(new_n466), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n472), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n481), .A2(G135), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n632), .A2(KEYINPUT80), .B1(G123), .B2(new_n483), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n633), .B(new_n635), .C1(KEYINPUT80), .C2(new_n632), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2435), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2438), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT14), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n644), .B(new_n649), .Z(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(G14), .ZN(G401));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n655), .B2(new_n652), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n673), .B2(KEYINPUT20), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(KEYINPUT20), .C2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  AND2_X1   g259(.A1(KEYINPUT24), .A2(G34), .ZN(new_n685));
  NOR2_X1   g260(.A1(KEYINPUT24), .A2(G34), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n685), .A2(new_n686), .A3(G29), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n479), .B2(G29), .ZN(new_n688));
  INV_X1    g263(.A(G2084), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT90), .Z(new_n691));
  NOR2_X1   g266(.A1(G29), .A2(G32), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n483), .A2(G129), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT89), .Z(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2090), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n705), .B(new_n706), .S(KEYINPUT91), .Z(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n704), .A2(G26), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n483), .A2(G128), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(G104), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n481), .A2(G140), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(G29), .ZN(new_n717));
  MUX2_X1   g292(.A(new_n709), .B(new_n717), .S(KEYINPUT28), .Z(new_n718));
  INV_X1    g293(.A(G2067), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n612), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G4), .B2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G1348), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n563), .B2(new_n721), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n707), .A2(new_n703), .B1(G1341), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n708), .A2(new_n720), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G1341), .B2(new_n728), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n688), .A2(new_n689), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(KEYINPUT30), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n636), .B2(new_n704), .ZN(new_n737));
  NOR2_X1   g312(.A1(G5), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G171), .B2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n737), .B1(G1961), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(G16), .A2(G21), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G286), .B2(new_n721), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n740), .B1(G1961), .B2(new_n739), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI211_X1 g319(.A(new_n733), .B(new_n744), .C1(new_n743), .C2(new_n742), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n626), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(new_n460), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT88), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G139), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n472), .A2(G103), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AND3_X1   g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G29), .B2(G33), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(G299), .A2(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT23), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n721), .A2(G20), .ZN(new_n760));
  MUX2_X1   g335(.A(KEYINPUT23), .B(new_n759), .S(new_n760), .Z(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(G1956), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n745), .A2(new_n756), .A3(new_n757), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(G1956), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n704), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n704), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n764), .B(new_n768), .C1(new_n754), .C2(new_n755), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n732), .A2(new_n763), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n721), .A2(G22), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G166), .B2(new_n721), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT86), .B(G1971), .Z(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n721), .A2(G6), .ZN(new_n775));
  INV_X1    g350(.A(G305), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n721), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT32), .B(G1981), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT85), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n777), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n772), .A2(new_n773), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n721), .A2(G23), .ZN(new_n782));
  INV_X1    g357(.A(G288), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n721), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1976), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n774), .A2(new_n780), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT34), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n481), .A2(G131), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n483), .A2(G119), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G24), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n602), .B(KEYINPUT84), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1986), .Z(new_n800));
  NAND3_X1  g375(.A1(new_n788), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT36), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n788), .A2(new_n803), .A3(new_n796), .A4(new_n800), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n691), .B(new_n770), .C1(new_n802), .C2(new_n804), .ZN(G311));
  AOI21_X1  g380(.A(new_n770), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  INV_X1    g381(.A(new_n691), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(G150));
  NAND2_X1  g383(.A1(new_n612), .A2(G559), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n620), .A2(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  INV_X1    g387(.A(G67), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n533), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G651), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT95), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n534), .A2(G93), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n526), .A2(G55), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n811), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT97), .B1(new_n563), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n620), .A2(KEYINPUT96), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n822), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n811), .B2(new_n819), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n810), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n832));
  OR3_X1    g407(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT39), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n832), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n819), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  XOR2_X1   g415(.A(new_n698), .B(KEYINPUT102), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n628), .B(new_n636), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n489), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n492), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT68), .B1(new_n492), .B2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n496), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n494), .A2(KEYINPUT69), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n849), .A2(new_n850), .B1(new_n501), .B2(new_n502), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n509), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n752), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n509), .A3(new_n851), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n479), .B(KEYINPUT99), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n487), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n483), .A2(G130), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT100), .Z(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  INV_X1    g437(.A(G118), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(G2105), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n460), .A2(KEYINPUT101), .A3(G118), .ZN(new_n865));
  OAI221_X1 g440(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G142), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n793), .ZN(new_n869));
  INV_X1    g444(.A(new_n716), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n857), .B(G162), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n853), .A3(new_n855), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n859), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n859), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n844), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n859), .A2(new_n873), .ZN(new_n878));
  INV_X1    g453(.A(new_n871), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n843), .A3(new_n874), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g459(.A(new_n828), .B(new_n623), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n612), .B(G299), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT41), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n602), .B(KEYINPUT103), .ZN(new_n893));
  NAND2_X1  g468(.A1(G303), .A2(new_n783), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n520), .B(G288), .C1(new_n536), .C2(new_n537), .ZN(new_n895));
  AOI21_X1  g470(.A(G305), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(G305), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  INV_X1    g475(.A(new_n893), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n900), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n890), .A2(new_n891), .ZN(new_n905));
  AND4_X1   g480(.A1(KEYINPUT104), .A2(new_n892), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n892), .A2(new_n905), .B1(KEYINPUT104), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n819), .A2(new_n604), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NOR2_X1   g487(.A1(G171), .A2(KEYINPUT105), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n825), .A2(new_n827), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n825), .B2(new_n827), .ZN(new_n917));
  AOI21_X1  g492(.A(G286), .B1(KEYINPUT105), .B2(G171), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n828), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n887), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n916), .B2(new_n917), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n918), .A3(new_n915), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n886), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n903), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n882), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n903), .B1(new_n926), .B2(new_n923), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n886), .B(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n934));
  OAI221_X1 g509(.A(new_n933), .B1(KEYINPUT106), .B2(new_n934), .C1(new_n920), .C2(new_n922), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n903), .B1(new_n935), .B2(new_n926), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n928), .A2(new_n936), .A3(KEYINPUT43), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n912), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n928), .ZN(new_n939));
  INV_X1    g514(.A(new_n929), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT43), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n928), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n944), .ZN(G397));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n852), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT107), .B(G40), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n469), .A2(new_n477), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n716), .B(new_n719), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT108), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n698), .B(G1996), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n793), .A2(new_n795), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n870), .A2(new_n719), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n954), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n954), .B1(new_n956), .B2(new_n698), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n954), .A2(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n793), .A2(new_n795), .ZN(new_n968));
  INV_X1    g543(.A(new_n959), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n958), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n953), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n953), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT48), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n962), .B(new_n967), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT63), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n584), .A2(G1976), .A3(new_n585), .A4(new_n586), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n509), .B2(new_n851), .ZN(new_n981));
  AOI211_X1 g556(.A(new_n978), .B(new_n980), .C1(new_n981), .C2(new_n951), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(KEYINPUT111), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n591), .A2(new_n593), .A3(new_n988), .A4(new_n595), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n542), .A2(G48), .A3(G543), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n990), .B(new_n592), .C1(new_n991), .C2(new_n515), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G1981), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT49), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT112), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n978), .B1(new_n981), .B2(new_n951), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n1001), .B(KEYINPUT49), .C1(new_n989), .C2(new_n993), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n997), .B(new_n998), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1004));
  AOI211_X1 g579(.A(new_n984), .B(new_n987), .C1(new_n999), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n513), .A2(new_n946), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n952), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  AND4_X1   g589(.A1(new_n1013), .A2(new_n852), .A3(new_n1014), .A4(new_n946), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1013), .B1(new_n981), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT110), .B(G2090), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n952), .B1(new_n1011), .B2(new_n948), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1971), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1010), .B(G8), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n513), .A2(new_n1014), .A3(new_n946), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n951), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1025), .A2(new_n1029), .A3(new_n1026), .A4(new_n951), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1019), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1023), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n978), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1005), .B(new_n1024), .C1(new_n1034), .C2(new_n1010), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(new_n952), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n743), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1012), .A2(new_n1017), .A3(new_n689), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n978), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G168), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n976), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1010), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n976), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1043), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1024), .A3(new_n1005), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1024), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1005), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n998), .B(KEYINPUT114), .Z(new_n1053));
  NAND2_X1  g628(.A1(new_n783), .A2(new_n985), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT115), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n999), .B2(new_n1004), .ZN(new_n1056));
  INV_X1    g631(.A(new_n989), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1038), .A2(new_n767), .A3(new_n949), .A4(new_n951), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1037), .A2(KEYINPUT123), .A3(new_n1038), .A4(new_n767), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT53), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1018), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1021), .A2(new_n767), .A3(new_n1022), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G286), .A2(G8), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT121), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1042), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1077), .B(KEYINPUT51), .C1(new_n1042), .C2(new_n1079), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1079), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1075), .A2(new_n1076), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1070), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT124), .B1(new_n1070), .B2(G171), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1014), .B1(new_n513), .B2(new_n946), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n1092), .A2(new_n1015), .A3(new_n1016), .A4(new_n952), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1093), .B2(G1961), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1068), .A2(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1022), .A2(G40), .A3(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n479), .A3(new_n1036), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1018), .A2(KEYINPUT125), .A3(new_n1065), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT54), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(KEYINPUT127), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT127), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1094), .A2(new_n1098), .A3(new_n1104), .A4(new_n1099), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(G171), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1070), .B2(G301), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1090), .A2(new_n1102), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1027), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1011), .A2(new_n948), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n951), .A3(new_n1022), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1018), .A2(new_n724), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n952), .A2(new_n947), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n719), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1116), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G299), .B(KEYINPUT57), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT117), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1111), .A2(new_n1114), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n612), .A2(new_n1122), .B1(new_n1127), .B2(KEYINPUT118), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1127), .A2(KEYINPUT118), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1117), .B(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  INV_X1    g707(.A(new_n612), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1121), .C1(new_n1093), .C2(G1348), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1348), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1121), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n612), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1119), .A2(new_n1132), .A3(new_n612), .A4(new_n1121), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1131), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(G1996), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT119), .B(G1341), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1120), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n563), .B(new_n1145), .C1(new_n1147), .C2(new_n1150), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1144), .A2(KEYINPUT59), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1130), .B1(new_n1143), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1087), .B1(new_n1109), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1075), .A2(KEYINPUT62), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1082), .A2(new_n1083), .B1(new_n1085), .B2(new_n1079), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1035), .A2(KEYINPUT126), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1035), .A2(KEYINPUT126), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1156), .A2(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1059), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n970), .B1(G1986), .B2(G290), .ZN(new_n1162));
  INV_X1    g737(.A(new_n972), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n954), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n975), .B1(new_n1161), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g740(.A1(new_n683), .A2(G319), .ZN(new_n1167));
  NOR2_X1   g741(.A1(G401), .A2(G227), .ZN(new_n1168));
  NAND2_X1  g742(.A1(new_n883), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g743(.A(new_n936), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n939), .A2(new_n1170), .A3(new_n942), .ZN(new_n1171));
  AOI211_X1 g745(.A(new_n1167), .B(new_n1169), .C1(new_n930), .C2(new_n1171), .ZN(G308));
  AOI21_X1  g746(.A(new_n1167), .B1(new_n1171), .B2(new_n930), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n1173), .A2(new_n883), .A3(new_n1168), .ZN(G225));
endmodule


