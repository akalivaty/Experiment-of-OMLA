//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n455), .A2(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n463), .B1(new_n475), .B2(new_n476), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(new_n475), .B2(new_n476), .ZN(new_n488));
  AND2_X1   g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n475), .B2(new_n476), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n463), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(G88), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n505), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n507), .A2(G89), .A3(new_n514), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n501), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n516), .A2(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n507), .A2(new_n514), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G171));
  AND2_X1   g108(.A1(new_n507), .A2(new_n514), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G81), .B1(G43), .B2(new_n516), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n504), .A2(new_n506), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n503), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n507), .A2(G91), .A3(new_n514), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n501), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n516), .A2(G53), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n513), .ZN(new_n558));
  OAI211_X1 g133(.A(G53), .B(G543), .C1(new_n558), .C2(new_n511), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT70), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n553), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NAND2_X1  g142(.A1(new_n525), .A2(KEYINPUT71), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n522), .A2(new_n524), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n569), .A2(new_n570), .A3(new_n520), .A4(new_n521), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  AOI22_X1  g148(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n515), .B(new_n517), .C1(new_n574), .C2(new_n501), .ZN(G303));
  OAI21_X1  g150(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n516), .A2(G49), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n530), .ZN(G288));
  NAND2_X1  g154(.A1(new_n516), .A2(G48), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n530), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n507), .A2(G61), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n501), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n516), .A2(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n530), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n507), .A2(G60), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n501), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT72), .B1(new_n590), .B2(new_n594), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(new_n514), .A2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT73), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G54), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n530), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT74), .B(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n539), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n602), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  MUX2_X1   g188(.A(G301), .B(new_n612), .S(new_n613), .Z(G284));
  MUX2_X1   g189(.A(G301), .B(new_n612), .S(new_n613), .Z(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n565), .B(KEYINPUT75), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  INV_X1    g194(.A(G860), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n612), .B1(G559), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT76), .ZN(G148));
  NOR2_X1   g197(.A1(new_n612), .A2(G559), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n544), .A2(new_n613), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT11), .Z(G282));
  INV_X1    g202(.A(new_n626), .ZN(G323));
  OR3_X1    g203(.A1(new_n478), .A2(KEYINPUT12), .A3(new_n474), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT12), .B1(new_n478), .B2(new_n474), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  MUX2_X1   g210(.A(G99), .B(G111), .S(G2105), .Z(new_n636));
  AOI22_X1  g211(.A1(G123), .A2(new_n481), .B1(new_n636), .B2(G2104), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n478), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT77), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT78), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT79), .Z(new_n661));
  NOR2_X1   g236(.A1(G2072), .A2(G2078), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n444), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(KEYINPUT17), .Z(new_n668));
  OAI211_X1 g243(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n661), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n661), .A3(new_n666), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n663), .A2(new_n660), .A3(new_n666), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT80), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2096), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT81), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G6), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n586), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G22), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G166), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(G16), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n704));
  NAND2_X1  g279(.A1(G288), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n534), .A2(G87), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n706), .A2(KEYINPUT85), .A3(new_n576), .A4(new_n577), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT33), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT86), .B(G1976), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n698), .B(new_n702), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n717));
  XNOR2_X1  g292(.A(G290), .B(KEYINPUT84), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G1986), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n709), .A2(G24), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT83), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n720), .B1(new_n719), .B2(new_n722), .ZN(new_n724));
  MUX2_X1   g299(.A(G95), .B(G107), .S(G2105), .Z(new_n725));
  AOI22_X1  g300(.A1(G119), .A2(new_n481), .B1(new_n725), .B2(G2104), .ZN(new_n726));
  INV_X1    g301(.A(G131), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n478), .ZN(new_n728));
  MUX2_X1   g303(.A(G25), .B(new_n728), .S(G29), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT82), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT87), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n716), .A2(new_n717), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G19), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n544), .B2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT89), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1341), .ZN(new_n740));
  NOR2_X1   g315(.A1(G4), .A2(G16), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT88), .Z(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n612), .B2(new_n709), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1348), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n749), .A2(G104), .A3(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G104), .ZN(new_n751));
  AOI21_X1  g326(.A(KEYINPUT90), .B1(new_n751), .B2(new_n463), .ZN(new_n752));
  OAI221_X1 g327(.A(G2104), .B1(G116), .B2(new_n463), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n481), .A2(G128), .ZN(new_n755));
  INV_X1    g330(.A(G140), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n478), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n748), .B1(new_n759), .B2(new_n746), .ZN(new_n760));
  INV_X1    g335(.A(G2067), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n744), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(KEYINPUT92), .B1(new_n740), .B2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G1341), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n739), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n762), .A4(new_n744), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n746), .A2(G35), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT101), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n746), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n764), .B(new_n768), .C1(G2090), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n709), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT102), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(G1956), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(G1956), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n772), .A2(G2090), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT103), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n716), .A2(KEYINPUT36), .A3(new_n717), .A4(new_n733), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n479), .A2(G139), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n785), .B(new_n788), .C1(new_n463), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(G164), .A2(G29), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G27), .B2(G29), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(new_n443), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n746), .A2(G32), .ZN(new_n797));
  NAND3_X1  g372(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT26), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n474), .A2(G2105), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(G105), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n479), .A2(G141), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n481), .A2(G129), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n797), .B1(new_n805), .B2(new_n746), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT27), .B(G1996), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n795), .A2(new_n443), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT31), .B(G11), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT30), .B(G28), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n746), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n639), .B2(new_n746), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n796), .A2(new_n809), .A3(new_n810), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G160), .A2(G29), .ZN(new_n817));
  AND2_X1   g392(.A1(KEYINPUT24), .A2(G34), .ZN(new_n818));
  NOR2_X1   g393(.A1(KEYINPUT24), .A2(G34), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n746), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G2084), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT95), .Z(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  NOR2_X1   g400(.A1(G171), .A2(new_n709), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G5), .B2(new_n709), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n793), .A2(new_n816), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n525), .A2(new_n709), .ZN(new_n831));
  MUX2_X1   g406(.A(new_n830), .B(KEYINPUT96), .S(new_n831), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1966), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n827), .A2(new_n825), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n806), .A2(new_n808), .B1(new_n822), .B2(new_n821), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n829), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND4_X1   g416(.A1(new_n736), .A2(new_n783), .A3(new_n784), .A4(new_n841), .ZN(G311));
  NAND4_X1  g417(.A1(new_n783), .A2(new_n736), .A3(new_n841), .A4(new_n784), .ZN(G150));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT104), .B(G55), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n530), .A2(new_n844), .B1(new_n600), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n507), .A2(G67), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n501), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n846), .B2(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  AND3_X1   g431(.A1(new_n602), .A2(new_n607), .A3(new_n611), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n851), .A2(new_n543), .A3(new_n853), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n543), .A2(new_n850), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n859), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(new_n620), .C1(new_n865), .C2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n856), .B1(new_n868), .B2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(new_n485), .B(G160), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n639), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n631), .B(new_n728), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n479), .A2(G142), .B1(G130), .B2(new_n481), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n463), .A2(KEYINPUT107), .A3(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT107), .B1(new_n463), .B2(G118), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n874), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT108), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n758), .B(G164), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n790), .B(new_n804), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(KEYINPUT109), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n886), .A2(KEYINPUT109), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n873), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT110), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n873), .A3(new_n886), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT40), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n896), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n899), .A2(new_n889), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n901), .ZN(G395));
  OR2_X1    g477(.A1(new_n862), .A2(new_n623), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n857), .A2(new_n565), .ZN(new_n904));
  NAND2_X1  g479(.A1(G299), .A2(new_n612), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n862), .A2(new_n623), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT41), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n903), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n862), .A2(new_n623), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(G290), .A2(new_n705), .A3(new_n707), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n708), .A2(new_n598), .A3(new_n597), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G166), .A2(KEYINPUT111), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  NAND2_X1  g496(.A1(G303), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n586), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(G305), .A3(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n917), .A2(new_n924), .A3(new_n925), .A4(new_n918), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT112), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n916), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n930), .A2(KEYINPUT112), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n911), .A2(new_n915), .A3(new_n929), .A4(new_n931), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n854), .A2(G868), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n938), .A2(KEYINPUT113), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT113), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  AND2_X1   g518(.A1(new_n938), .A2(new_n940), .ZN(G331));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g520(.A1(G301), .A2(G168), .ZN(new_n946));
  NAND3_X1  g521(.A1(G171), .A2(new_n568), .A3(new_n571), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n862), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n860), .A2(new_n861), .A3(new_n946), .A4(new_n947), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT114), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n862), .A2(new_n952), .A3(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n908), .A2(new_n910), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n950), .ZN(new_n956));
  OAI22_X1  g531(.A1(new_n954), .A2(new_n955), .B1(new_n906), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n927), .B2(new_n928), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n927), .A2(new_n958), .A3(new_n928), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n954), .A2(new_n912), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n908), .A3(new_n910), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n929), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n896), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(new_n963), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n906), .B1(new_n951), .B2(new_n953), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n967), .A2(new_n968), .B1(new_n960), .B2(new_n959), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n964), .A3(new_n970), .A4(new_n896), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n945), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n964), .A3(new_n896), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT43), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n961), .A2(new_n970), .A3(new_n896), .A4(new_n964), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n973), .B2(KEYINPUT43), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n972), .B1(new_n979), .B2(new_n945), .ZN(G397));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n499), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G160), .A2(G40), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n758), .B(new_n761), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n804), .B(G1996), .Z(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n728), .A2(new_n731), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n990), .A2(new_n991), .B1(G2067), .B2(new_n758), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n986), .B1(new_n992), .B2(KEYINPUT127), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n986), .A2(new_n720), .A3(new_n598), .A4(new_n597), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT48), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(new_n988), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n728), .B(new_n731), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n986), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT48), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n995), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n993), .A2(new_n994), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n987), .B1(new_n988), .B2(new_n805), .ZN(new_n1004));
  OR3_X1    g579(.A1(new_n987), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT46), .B1(new_n987), .B2(G1996), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT47), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n525), .A2(KEYINPUT122), .A3(G8), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT122), .B1(new_n525), .B2(G8), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n1012), .B2(KEYINPUT124), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n982), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n981), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n985), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1019));
  INV_X1    g594(.A(G40), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n468), .A2(new_n471), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n984), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n822), .A2(new_n1018), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1012), .B(new_n1014), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT51), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(KEYINPUT4), .A2(G138), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n464), .B2(new_n465), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n493), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1032), .A2(new_n463), .B1(new_n497), .B2(new_n496), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n1033), .B2(new_n490), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1021), .B1(new_n1034), .B2(KEYINPUT45), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1019), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1023), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n981), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT50), .B1(new_n499), .B2(new_n981), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n822), .B(new_n1021), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1025), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1029), .B1(new_n1041), .B2(new_n1027), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT123), .B1(new_n1043), .B2(new_n1027), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n1045), .B(new_n1012), .C1(new_n1037), .C2(new_n1040), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1026), .B(new_n1042), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(KEYINPUT123), .A3(new_n1027), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(KEYINPUT62), .A3(new_n1026), .A4(new_n1042), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2090), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1059), .A2(new_n1018), .B1(new_n1022), .B2(new_n701), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n1025), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1021), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1063));
  OAI22_X1  g638(.A1(new_n1062), .A2(G1971), .B1(new_n1063), .B2(G2090), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1058), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(G8), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n982), .A2(new_n985), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n1025), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n705), .A2(new_n707), .A3(G1976), .ZN(new_n1069));
  INV_X1    g644(.A(G1976), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(G288), .B2(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1034), .A2(new_n1021), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(new_n582), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n583), .A2(new_n584), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G651), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(G1981), .B1(new_n582), .B2(new_n585), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT49), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1061), .A2(new_n1066), .A3(new_n1075), .A4(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n984), .A2(new_n443), .A3(new_n1019), .A4(new_n1021), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1063), .A2(new_n825), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(G2078), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n984), .A2(new_n1019), .A3(new_n1021), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1092), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1054), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1060), .A2(new_n1025), .A3(new_n1058), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n1091), .A3(new_n1075), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G288), .A2(G1976), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1091), .A2(new_n1105), .B1(new_n1079), .B2(new_n586), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1106), .B2(new_n1077), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1041), .A2(new_n1109), .A3(new_n572), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1041), .B2(new_n572), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1108), .B1(new_n1112), .B2(new_n1092), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1041), .A2(new_n572), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1041), .A2(new_n1109), .A3(new_n572), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1065), .B1(new_n1064), .B2(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1103), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1075), .A2(new_n1091), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(KEYINPUT63), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1107), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1063), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1067), .A2(new_n761), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n612), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g702(.A(new_n561), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n553), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT120), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(new_n1127), .C1(new_n553), .C2(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n562), .A2(new_n564), .ZN(new_n1133));
  INV_X1    g708(.A(new_n553), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT57), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G1956), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1063), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT56), .B(G2072), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n984), .A2(new_n1019), .A3(new_n1021), .A4(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1126), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1141), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1124), .A2(new_n612), .A3(new_n1125), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT60), .B1(new_n1151), .B2(new_n1126), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n612), .A2(KEYINPUT60), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1124), .A2(new_n1125), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1145), .A2(KEYINPUT61), .A3(new_n1141), .ZN(new_n1155));
  AND4_X1   g730(.A1(new_n1150), .A2(new_n1152), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT58), .B(G1341), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1022), .A2(G1996), .B1(new_n1067), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(KEYINPUT121), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1158), .A2(KEYINPUT121), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n544), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT59), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n544), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1146), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1095), .A2(new_n1096), .A3(G301), .A4(new_n1098), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1100), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT54), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1100), .A2(KEYINPUT54), .A3(new_n1167), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1092), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1173), .A2(new_n1175), .A3(new_n1047), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1102), .B(new_n1122), .C1(new_n1166), .C2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(G290), .B(new_n720), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1000), .B1(new_n987), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT117), .Z(new_n1180));
  AND3_X1   g755(.A1(new_n1177), .A2(KEYINPUT126), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT126), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1009), .B1(new_n1181), .B2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g758(.A1(G227), .A2(new_n461), .A3(G401), .A4(G229), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n889), .B2(new_n899), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n979), .A2(new_n1186), .ZN(G308));
  OAI221_X1 g761(.A(new_n1185), .B1(new_n889), .B2(new_n899), .C1(new_n977), .C2(new_n978), .ZN(G225));
endmodule


