

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754;

  XNOR2_X1 U368 ( .A(n408), .B(KEYINPUT32), .ZN(n752) );
  OR2_X1 U369 ( .A1(n574), .A2(n406), .ZN(n408) );
  NOR2_X1 U370 ( .A1(n671), .A2(n672), .ZN(n559) );
  XNOR2_X1 U371 ( .A(n490), .B(n350), .ZN(n671) );
  NOR2_X1 U372 ( .A1(n632), .A2(G902), .ZN(n443) );
  XNOR2_X1 U373 ( .A(n459), .B(n489), .ZN(n350) );
  XNOR2_X1 U374 ( .A(n410), .B(n734), .ZN(n705) );
  XNOR2_X1 U375 ( .A(n511), .B(n347), .ZN(n734) );
  XNOR2_X1 U376 ( .A(n349), .B(n355), .ZN(n482) );
  XNOR2_X1 U377 ( .A(n481), .B(KEYINPUT74), .ZN(n349) );
  XNOR2_X1 U378 ( .A(KEYINPUT16), .B(G122), .ZN(n347) );
  BUF_X1 U379 ( .A(G113), .Z(n348) );
  INV_X2 U380 ( .A(G953), .ZN(n733) );
  AND2_X2 U381 ( .A1(n645), .A2(n752), .ZN(n553) );
  NAND2_X2 U382 ( .A1(n456), .A2(n365), .ZN(n398) );
  INV_X2 U383 ( .A(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U384 ( .A(G116), .B(G113), .ZN(n458) );
  NOR2_X2 U385 ( .A1(n712), .A2(G902), .ZN(n490) );
  XNOR2_X2 U386 ( .A(n603), .B(KEYINPUT41), .ZN(n692) );
  NOR2_X2 U387 ( .A1(n693), .A2(n564), .ZN(n515) );
  XNOR2_X2 U388 ( .A(n403), .B(n514), .ZN(n693) );
  AND2_X2 U389 ( .A1(n396), .A2(n395), .ZN(n394) );
  NOR2_X2 U390 ( .A1(n663), .A2(n664), .ZN(n603) );
  XNOR2_X2 U391 ( .A(n584), .B(KEYINPUT39), .ZN(n605) );
  NAND2_X1 U392 ( .A1(n394), .A2(n391), .ZN(n730) );
  NOR2_X1 U393 ( .A1(n588), .A2(n586), .ZN(n561) );
  INV_X1 U394 ( .A(G217), .ZN(n452) );
  NAND2_X1 U395 ( .A1(n393), .A2(n358), .ZN(n391) );
  AND2_X1 U396 ( .A1(n573), .A2(n392), .ZN(n358) );
  NOR2_X1 U397 ( .A1(n750), .A2(n754), .ZN(n418) );
  XNOR2_X1 U398 ( .A(n606), .B(n409), .ZN(n750) );
  XNOR2_X1 U399 ( .A(n548), .B(n547), .ZN(n574) );
  XNOR2_X1 U400 ( .A(n604), .B(KEYINPUT42), .ZN(n754) );
  INV_X1 U401 ( .A(n599), .ZN(n678) );
  XNOR2_X1 U402 ( .A(n715), .B(n460), .ZN(n716) );
  XNOR2_X1 U403 ( .A(n405), .B(G125), .ZN(n379) );
  XNOR2_X1 U404 ( .A(KEYINPUT75), .B(G101), .ZN(n462) );
  INV_X1 U405 ( .A(G146), .ZN(n405) );
  XNOR2_X1 U406 ( .A(n457), .B(n463), .ZN(n511) );
  XNOR2_X1 U407 ( .A(n462), .B(n458), .ZN(n457) );
  BUF_X1 U408 ( .A(n730), .Z(n351) );
  XNOR2_X1 U409 ( .A(n490), .B(n489), .ZN(n352) );
  BUF_X1 U410 ( .A(n559), .Z(n353) );
  XNOR2_X2 U411 ( .A(n742), .B(G146), .ZN(n513) );
  XNOR2_X2 U412 ( .A(n482), .B(n483), .ZN(n742) );
  INV_X1 U413 ( .A(n657), .ZN(n437) );
  NAND2_X1 U414 ( .A1(n556), .A2(n544), .ZN(n663) );
  NAND2_X1 U415 ( .A1(n450), .A2(n389), .ZN(n376) );
  NOR2_X1 U416 ( .A1(n404), .A2(n572), .ZN(n389) );
  XOR2_X1 U417 ( .A(G140), .B(KEYINPUT73), .Z(n493) );
  NOR2_X1 U418 ( .A1(n390), .A2(n376), .ZN(n393) );
  INV_X1 U419 ( .A(n398), .ZN(n390) );
  XNOR2_X1 U420 ( .A(n442), .B(G128), .ZN(n480) );
  INV_X1 U421 ( .A(G143), .ZN(n442) );
  XOR2_X1 U422 ( .A(KEYINPUT90), .B(KEYINPUT17), .Z(n467) );
  XNOR2_X1 U423 ( .A(n440), .B(n439), .ZN(n664) );
  INV_X1 U424 ( .A(KEYINPUT111), .ZN(n439) );
  NAND2_X1 U425 ( .A1(n661), .A2(n660), .ZN(n440) );
  INV_X1 U426 ( .A(KEYINPUT77), .ZN(n373) );
  NAND2_X1 U427 ( .A1(n375), .A2(KEYINPUT77), .ZN(n374) );
  NAND2_X1 U428 ( .A1(n580), .A2(n373), .ZN(n369) );
  NOR2_X1 U429 ( .A1(n361), .A2(n448), .ZN(n447) );
  INV_X1 U430 ( .A(n753), .ZN(n448) );
  XNOR2_X1 U431 ( .A(n480), .B(n441), .ZN(n521) );
  INV_X1 U432 ( .A(G134), .ZN(n441) );
  XNOR2_X1 U433 ( .A(G116), .B(G122), .ZN(n516) );
  XOR2_X1 U434 ( .A(KEYINPUT9), .B(G107), .Z(n517) );
  XNOR2_X1 U435 ( .A(n423), .B(n422), .ZN(n591) );
  INV_X1 U436 ( .A(KEYINPUT104), .ZN(n422) );
  NAND2_X1 U437 ( .A1(n424), .A2(n651), .ZN(n423) );
  INV_X1 U438 ( .A(n623), .ZN(n428) );
  XNOR2_X1 U439 ( .A(n402), .B(n401), .ZN(n609) );
  INV_X1 U440 ( .A(KEYINPUT19), .ZN(n401) );
  XNOR2_X1 U441 ( .A(n537), .B(n400), .ZN(n557) );
  XNOR2_X1 U442 ( .A(n538), .B(G475), .ZN(n400) );
  NOR2_X1 U443 ( .A1(n720), .A2(G902), .ZN(n523) );
  XNOR2_X1 U444 ( .A(n546), .B(KEYINPUT67), .ZN(n547) );
  NAND2_X1 U445 ( .A1(n415), .A2(n359), .ZN(n548) );
  XNOR2_X1 U446 ( .A(n366), .B(n492), .ZN(n505) );
  NOR2_X1 U447 ( .A1(G952), .A2(n733), .ZN(n724) );
  XNOR2_X1 U448 ( .A(n607), .B(n608), .ZN(n409) );
  NAND2_X1 U449 ( .A1(KEYINPUT44), .A2(n382), .ZN(n381) );
  INV_X1 U450 ( .A(KEYINPUT87), .ZN(n382) );
  OR2_X1 U451 ( .A1(G237), .A2(G902), .ZN(n470) );
  XNOR2_X1 U452 ( .A(n367), .B(KEYINPUT20), .ZN(n506) );
  NAND2_X1 U453 ( .A1(n491), .A2(G234), .ZN(n367) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n413) );
  XOR2_X1 U455 ( .A(KEYINPUT89), .B(n461), .Z(n629) );
  XNOR2_X1 U456 ( .A(n368), .B(KEYINPUT15), .ZN(n461) );
  INV_X1 U457 ( .A(G902), .ZN(n368) );
  XNOR2_X1 U458 ( .A(n493), .B(n354), .ZN(n484) );
  NAND2_X1 U459 ( .A1(G234), .A2(G237), .ZN(n472) );
  AND2_X1 U460 ( .A1(n590), .A2(n425), .ZN(n424) );
  INV_X1 U461 ( .A(n598), .ZN(n425) );
  NAND2_X1 U462 ( .A1(n506), .A2(G217), .ZN(n366) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n509) );
  XNOR2_X1 U464 ( .A(n421), .B(n420), .ZN(n735) );
  INV_X1 U465 ( .A(G110), .ZN(n420) );
  XNOR2_X1 U466 ( .A(G107), .B(G104), .ZN(n421) );
  XOR2_X1 U467 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n528) );
  XNOR2_X1 U468 ( .A(G131), .B(G140), .ZN(n527) );
  XNOR2_X1 U469 ( .A(n348), .B(G143), .ZN(n531) );
  XOR2_X1 U470 ( .A(G104), .B(G122), .Z(n532) );
  XOR2_X1 U471 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n526) );
  XNOR2_X1 U472 ( .A(n735), .B(KEYINPUT76), .ZN(n485) );
  INV_X1 U473 ( .A(n480), .ZN(n434) );
  XNOR2_X1 U474 ( .A(n356), .B(n379), .ZN(n465) );
  XNOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT18), .ZN(n466) );
  AND2_X1 U476 ( .A1(n370), .A2(n357), .ZN(n622) );
  NAND2_X1 U477 ( .A1(n587), .A2(n373), .ZN(n372) );
  INV_X1 U478 ( .A(KEYINPUT93), .ZN(n562) );
  INV_X1 U479 ( .A(KEYINPUT0), .ZN(n478) );
  XNOR2_X1 U480 ( .A(n632), .B(KEYINPUT62), .ZN(n633) );
  INV_X1 U481 ( .A(n745), .ZN(n383) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n720) );
  XNOR2_X1 U483 ( .A(n520), .B(n362), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n521), .B(n519), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n696), .B(n417), .ZN(n416) );
  INV_X1 U486 ( .A(KEYINPUT82), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n429) );
  AND2_X1 U488 ( .A1(n592), .A2(n412), .ZN(n431) );
  NAND2_X1 U489 ( .A1(n385), .A2(n597), .ZN(n657) );
  XNOR2_X1 U490 ( .A(n386), .B(n596), .ZN(n385) );
  NOR2_X1 U491 ( .A1(n594), .A2(n428), .ZN(n386) );
  NAND2_X1 U492 ( .A1(n549), .A2(n407), .ZN(n406) );
  XNOR2_X1 U493 ( .A(n558), .B(KEYINPUT101), .ZN(n651) );
  NOR2_X1 U494 ( .A1(n588), .A2(n575), .ZN(n638) );
  XNOR2_X1 U495 ( .A(n377), .B(KEYINPUT86), .ZN(n575) );
  NAND2_X1 U496 ( .A1(n412), .A2(n407), .ZN(n378) );
  AND2_X1 U497 ( .A1(n454), .A2(n725), .ZN(n726) );
  XNOR2_X1 U498 ( .A(n710), .B(n411), .ZN(n714) );
  XNOR2_X1 U499 ( .A(n713), .B(n711), .ZN(n411) );
  BUF_X1 U500 ( .A(n671), .Z(n412) );
  AND2_X1 U501 ( .A1(G227), .A2(n733), .ZN(n354) );
  XNOR2_X1 U502 ( .A(G131), .B(G137), .ZN(n355) );
  AND2_X1 U503 ( .A1(G224), .A2(n733), .ZN(n356) );
  AND2_X1 U504 ( .A1(n369), .A2(n372), .ZN(n357) );
  XNOR2_X1 U505 ( .A(KEYINPUT102), .B(n545), .ZN(n359) );
  XOR2_X1 U506 ( .A(G472), .B(KEYINPUT95), .Z(n360) );
  AND2_X1 U507 ( .A1(n429), .A2(n428), .ZN(n361) );
  XNOR2_X1 U508 ( .A(KEYINPUT99), .B(KEYINPUT7), .ZN(n362) );
  INV_X1 U509 ( .A(n590), .ZN(n407) );
  XOR2_X1 U510 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n363) );
  XOR2_X1 U511 ( .A(n723), .B(KEYINPUT122), .Z(n364) );
  AND2_X1 U512 ( .A1(KEYINPUT44), .A2(n543), .ZN(n365) );
  NOR2_X1 U513 ( .A1(n581), .A2(n371), .ZN(n370) );
  NOR2_X1 U514 ( .A1(n580), .A2(n374), .ZN(n371) );
  XNOR2_X2 U515 ( .A(n563), .B(n562), .ZN(n580) );
  INV_X1 U516 ( .A(n587), .ZN(n375) );
  NAND2_X1 U517 ( .A1(n376), .A2(n363), .ZN(n395) );
  OR2_X1 U518 ( .A1(n574), .A2(n378), .ZN(n377) );
  INV_X1 U519 ( .A(n379), .ZN(n380) );
  XNOR2_X1 U520 ( .A(n380), .B(KEYINPUT10), .ZN(n534) );
  NOR2_X1 U521 ( .A1(n419), .A2(n381), .ZN(n404) );
  XNOR2_X2 U522 ( .A(n542), .B(n541), .ZN(n419) );
  NOR2_X2 U523 ( .A1(n730), .A2(n384), .ZN(n630) );
  XNOR2_X1 U524 ( .A(n384), .B(n383), .ZN(n743) );
  NAND2_X1 U525 ( .A1(n449), .A2(n447), .ZN(n384) );
  XNOR2_X2 U526 ( .A(n388), .B(KEYINPUT71), .ZN(n481) );
  INV_X1 U527 ( .A(n363), .ZN(n392) );
  NAND2_X1 U528 ( .A1(n397), .A2(n363), .ZN(n396) );
  NAND2_X1 U529 ( .A1(n573), .A2(n398), .ZN(n397) );
  XNOR2_X1 U530 ( .A(n599), .B(KEYINPUT6), .ZN(n590) );
  NAND2_X1 U531 ( .A1(n552), .A2(n588), .ZN(n645) );
  XNOR2_X1 U532 ( .A(n399), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U533 ( .A1(n718), .A2(n724), .ZN(n399) );
  XNOR2_X1 U534 ( .A(n706), .B(n707), .ZN(n708) );
  NAND2_X1 U535 ( .A1(n722), .A2(G210), .ZN(n706) );
  NOR2_X4 U536 ( .A1(n631), .A2(n696), .ZN(n722) );
  NAND2_X2 U537 ( .A1(n630), .A2(KEYINPUT2), .ZN(n697) );
  NAND2_X1 U538 ( .A1(n471), .A2(n660), .ZN(n402) );
  NOR2_X1 U539 ( .A1(n437), .A2(n628), .ZN(n436) );
  NAND2_X1 U540 ( .A1(n559), .A2(n590), .ZN(n403) );
  NOR2_X1 U541 ( .A1(n723), .A2(G902), .ZN(n504) );
  NAND2_X1 U542 ( .A1(n438), .A2(n436), .ZN(n414) );
  XNOR2_X1 U543 ( .A(n414), .B(n413), .ZN(n449) );
  XNOR2_X1 U544 ( .A(n432), .B(n485), .ZN(n410) );
  INV_X1 U545 ( .A(n564), .ZN(n415) );
  XNOR2_X2 U546 ( .A(n479), .B(n478), .ZN(n564) );
  NOR2_X2 U547 ( .A1(n630), .A2(KEYINPUT2), .ZN(n696) );
  NOR2_X1 U548 ( .A1(n700), .A2(G953), .ZN(n701) );
  NAND2_X1 U549 ( .A1(n416), .A2(n697), .ZN(n698) );
  XNOR2_X1 U550 ( .A(n418), .B(KEYINPUT46), .ZN(n438) );
  NAND2_X1 U551 ( .A1(n419), .A2(KEYINPUT87), .ZN(n569) );
  XNOR2_X1 U552 ( .A(n419), .B(n751), .ZN(G24) );
  XNOR2_X1 U553 ( .A(n419), .B(n446), .ZN(n445) );
  XNOR2_X1 U554 ( .A(n593), .B(KEYINPUT107), .ZN(n430) );
  XNOR2_X1 U555 ( .A(n435), .B(n433), .ZN(n432) );
  XNOR2_X1 U556 ( .A(n481), .B(n434), .ZN(n433) );
  XNOR2_X1 U557 ( .A(n465), .B(n468), .ZN(n435) );
  INV_X1 U558 ( .A(n595), .ZN(n623) );
  XNOR2_X1 U559 ( .A(n595), .B(KEYINPUT38), .ZN(n661) );
  NAND2_X1 U560 ( .A1(n453), .A2(n451), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n455), .B(n364), .ZN(n454) );
  NAND2_X2 U562 ( .A1(n697), .A2(n629), .ZN(n631) );
  XNOR2_X2 U563 ( .A(n443), .B(n360), .ZN(n599) );
  XNOR2_X1 U564 ( .A(n513), .B(n512), .ZN(n632) );
  NAND2_X1 U565 ( .A1(n444), .A2(n543), .ZN(n554) );
  NAND2_X1 U566 ( .A1(n445), .A2(n571), .ZN(n444) );
  INV_X1 U567 ( .A(KEYINPUT69), .ZN(n446) );
  INV_X1 U568 ( .A(n638), .ZN(n450) );
  NOR2_X1 U569 ( .A1(n696), .A2(n452), .ZN(n451) );
  INV_X1 U570 ( .A(n631), .ZN(n453) );
  NAND2_X1 U571 ( .A1(n553), .A2(n446), .ZN(n456) );
  INV_X1 U572 ( .A(n588), .ZN(n674) );
  NOR2_X2 U573 ( .A1(n708), .A2(n724), .ZN(n709) );
  XOR2_X1 U574 ( .A(KEYINPUT68), .B(KEYINPUT1), .Z(n459) );
  XNOR2_X1 U575 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n460) );
  XNOR2_X1 U576 ( .A(KEYINPUT103), .B(KEYINPUT33), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U579 ( .A(n724), .ZN(n725) );
  XNOR2_X1 U580 ( .A(n717), .B(n716), .ZN(n718) );
  INV_X1 U581 ( .A(KEYINPUT109), .ZN(n608) );
  INV_X1 U582 ( .A(KEYINPUT63), .ZN(n636) );
  INV_X1 U583 ( .A(KEYINPUT65), .ZN(n543) );
  XOR2_X1 U584 ( .A(G119), .B(KEYINPUT3), .Z(n463) );
  XNOR2_X1 U585 ( .A(n467), .B(n466), .ZN(n468) );
  INV_X1 U586 ( .A(n629), .ZN(n491) );
  NAND2_X1 U587 ( .A1(n705), .A2(n491), .ZN(n583) );
  NAND2_X1 U588 ( .A1(G210), .A2(n470), .ZN(n582) );
  INV_X1 U589 ( .A(n582), .ZN(n469) );
  XNOR2_X1 U590 ( .A(n583), .B(n469), .ZN(n471) );
  NAND2_X1 U591 ( .A1(G214), .A2(n470), .ZN(n660) );
  XOR2_X1 U592 ( .A(KEYINPUT14), .B(KEYINPUT92), .Z(n473) );
  XOR2_X1 U593 ( .A(n473), .B(n472), .Z(n474) );
  NAND2_X1 U594 ( .A1(G952), .A2(n474), .ZN(n691) );
  NOR2_X1 U595 ( .A1(G953), .A2(n691), .ZN(n579) );
  AND2_X1 U596 ( .A1(n474), .A2(G953), .ZN(n475) );
  NAND2_X1 U597 ( .A1(G902), .A2(n475), .ZN(n577) );
  NOR2_X1 U598 ( .A1(G898), .A2(n577), .ZN(n476) );
  NOR2_X1 U599 ( .A1(n579), .A2(n476), .ZN(n477) );
  NOR2_X2 U600 ( .A1(n609), .A2(n477), .ZN(n479) );
  INV_X1 U601 ( .A(n521), .ZN(n483) );
  XNOR2_X1 U602 ( .A(G101), .B(KEYINPUT80), .ZN(n487) );
  XNOR2_X1 U603 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n513), .B(n488), .ZN(n712) );
  INV_X1 U605 ( .A(G469), .ZN(n489) );
  XOR2_X1 U606 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n492) );
  XOR2_X1 U607 ( .A(n493), .B(n534), .Z(n740) );
  XNOR2_X1 U608 ( .A(G119), .B(G137), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(KEYINPUT79), .ZN(n498) );
  XOR2_X1 U610 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n496) );
  XNOR2_X1 U611 ( .A(G128), .B(G110), .ZN(n495) );
  XNOR2_X1 U612 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U613 ( .A(n498), .B(n497), .Z(n502) );
  XOR2_X1 U614 ( .A(KEYINPUT72), .B(KEYINPUT8), .Z(n500) );
  NAND2_X1 U615 ( .A1(G234), .A2(n733), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n500), .B(n499), .ZN(n518) );
  NAND2_X1 U617 ( .A1(G221), .A2(n518), .ZN(n501) );
  XNOR2_X1 U618 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U619 ( .A(n740), .B(n503), .ZN(n723) );
  XNOR2_X2 U620 ( .A(n505), .B(n504), .ZN(n588) );
  NAND2_X1 U621 ( .A1(n506), .A2(G221), .ZN(n507) );
  XOR2_X1 U622 ( .A(n507), .B(KEYINPUT21), .Z(n675) );
  INV_X1 U623 ( .A(n675), .ZN(n586) );
  INV_X1 U624 ( .A(n561), .ZN(n672) );
  NOR2_X1 U625 ( .A1(G953), .A2(G237), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n524), .A2(G210), .ZN(n508) );
  XNOR2_X1 U627 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U628 ( .A(n515), .B(KEYINPUT34), .ZN(n539) );
  XNOR2_X1 U629 ( .A(n517), .B(n516), .ZN(n520) );
  NAND2_X1 U630 ( .A1(G217), .A2(n518), .ZN(n519) );
  XNOR2_X1 U631 ( .A(KEYINPUT100), .B(G478), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n523), .B(n522), .ZN(n556) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n538) );
  NAND2_X1 U634 ( .A1(G214), .A2(n524), .ZN(n525) );
  XNOR2_X1 U635 ( .A(n526), .B(n525), .ZN(n530) );
  XNOR2_X1 U636 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U637 ( .A(n530), .B(n529), .Z(n536) );
  XNOR2_X1 U638 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U639 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U640 ( .A(n536), .B(n535), .ZN(n715) );
  NOR2_X1 U641 ( .A1(G902), .A2(n715), .ZN(n537) );
  INV_X1 U642 ( .A(n557), .ZN(n544) );
  NOR2_X1 U643 ( .A1(n556), .A2(n544), .ZN(n625) );
  NAND2_X1 U644 ( .A1(n539), .A2(n625), .ZN(n542) );
  XOR2_X1 U645 ( .A(KEYINPUT35), .B(KEYINPUT85), .Z(n540) );
  XNOR2_X1 U646 ( .A(KEYINPUT81), .B(n540), .ZN(n541) );
  INV_X1 U647 ( .A(KEYINPUT44), .ZN(n571) );
  NOR2_X1 U648 ( .A1(n586), .A2(n663), .ZN(n545) );
  INV_X1 U649 ( .A(KEYINPUT22), .ZN(n546) );
  NOR2_X1 U650 ( .A1(n412), .A2(n674), .ZN(n549) );
  INV_X1 U651 ( .A(n412), .ZN(n597) );
  OR2_X1 U652 ( .A1(n597), .A2(n678), .ZN(n550) );
  NOR2_X1 U653 ( .A1(n574), .A2(n550), .ZN(n551) );
  XNOR2_X1 U654 ( .A(n551), .B(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n554), .A2(n553), .ZN(n573) );
  NOR2_X1 U656 ( .A1(KEYINPUT65), .A2(KEYINPUT87), .ZN(n555) );
  NOR2_X1 U657 ( .A1(KEYINPUT44), .A2(n555), .ZN(n568) );
  NOR2_X1 U658 ( .A1(n556), .A2(n557), .ZN(n653) );
  NAND2_X1 U659 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U660 ( .A1(n653), .A2(n651), .ZN(n665) );
  NAND2_X1 U661 ( .A1(n678), .A2(n353), .ZN(n682) );
  NOR2_X1 U662 ( .A1(n564), .A2(n682), .ZN(n560) );
  XOR2_X1 U663 ( .A(KEYINPUT31), .B(n560), .Z(n654) );
  NAND2_X1 U664 ( .A1(n561), .A2(n352), .ZN(n563) );
  OR2_X1 U665 ( .A1(n580), .A2(n564), .ZN(n565) );
  NOR2_X1 U666 ( .A1(n678), .A2(n565), .ZN(n641) );
  NOR2_X1 U667 ( .A1(n654), .A2(n641), .ZN(n566) );
  NOR2_X1 U668 ( .A1(n665), .A2(n566), .ZN(n567) );
  NOR2_X1 U669 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U671 ( .A1(n678), .A2(n660), .ZN(n576) );
  XNOR2_X1 U672 ( .A(KEYINPUT30), .B(n576), .ZN(n581) );
  NOR2_X1 U673 ( .A1(G900), .A2(n577), .ZN(n578) );
  NOR2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n587) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n622), .A2(n661), .ZN(n584) );
  NAND2_X1 U677 ( .A1(n653), .A2(n605), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n585), .B(KEYINPUT112), .ZN(n753) );
  NOR2_X1 U679 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n591), .A2(n660), .ZN(n594) );
  XNOR2_X1 U682 ( .A(n594), .B(KEYINPUT105), .ZN(n592) );
  XNOR2_X1 U683 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n593) );
  XNOR2_X1 U684 ( .A(KEYINPUT36), .B(KEYINPUT88), .ZN(n596) );
  NOR2_X1 U685 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U686 ( .A(KEYINPUT28), .B(n600), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n602), .A2(n352), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n610), .A2(n692), .ZN(n604) );
  XOR2_X1 U689 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n607) );
  NAND2_X1 U690 ( .A1(n605), .A2(n651), .ZN(n606) );
  NOR2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n649) );
  NOR2_X1 U692 ( .A1(n665), .A2(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U693 ( .A1(KEYINPUT70), .A2(n611), .ZN(n612) );
  NAND2_X1 U694 ( .A1(KEYINPUT84), .A2(n612), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n649), .A2(n613), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n649), .A2(KEYINPUT70), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n614), .A2(KEYINPUT84), .ZN(n616) );
  INV_X1 U698 ( .A(n665), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U700 ( .A1(KEYINPUT47), .A2(n617), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U702 ( .A1(KEYINPUT84), .A2(KEYINPUT47), .ZN(n620) );
  NOR2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n627) );
  AND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U705 ( .A(KEYINPUT108), .B(n624), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n648) );
  NAND2_X1 U707 ( .A1(n627), .A2(n648), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n722), .A2(G472), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X2 U710 ( .A1(n635), .A2(n724), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(n636), .ZN(G57) );
  XOR2_X1 U712 ( .A(n638), .B(G101), .Z(G3) );
  XOR2_X1 U713 ( .A(G104), .B(KEYINPUT113), .Z(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n651), .ZN(n639) );
  XNOR2_X1 U715 ( .A(n640), .B(n639), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n643) );
  NAND2_X1 U717 ( .A1(n641), .A2(n653), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U719 ( .A(G107), .B(n644), .ZN(G9) );
  XNOR2_X1 U720 ( .A(n645), .B(G110), .ZN(G12) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n647) );
  NAND2_X1 U722 ( .A1(n649), .A2(n653), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(G30) );
  XNOR2_X1 U724 ( .A(G143), .B(n648), .ZN(G45) );
  NAND2_X1 U725 ( .A1(n649), .A2(n651), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(G146), .ZN(G48) );
  NAND2_X1 U727 ( .A1(n654), .A2(n651), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(n348), .ZN(G15) );
  NAND2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(KEYINPUT114), .ZN(n656) );
  XNOR2_X1 U731 ( .A(G116), .B(n656), .ZN(G18) );
  XNOR2_X1 U732 ( .A(KEYINPUT37), .B(KEYINPUT115), .ZN(n658) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U734 ( .A(G125), .B(n659), .ZN(G27) );
  XOR2_X1 U735 ( .A(G140), .B(n361), .Z(G42) );
  NOR2_X1 U736 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n668) );
  NOR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n666), .B(KEYINPUT118), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n669), .A2(n693), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT119), .B(n670), .Z(n688) );
  NAND2_X1 U743 ( .A1(n672), .A2(n412), .ZN(n673) );
  XNOR2_X1 U744 ( .A(KEYINPUT50), .B(n673), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT49), .B(n676), .Z(n677) );
  NOR2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT116), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n685) );
  XOR2_X1 U751 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n686), .A2(n692), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U755 ( .A(n689), .B(KEYINPUT52), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n699) );
  NAND2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n701), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U761 ( .A(KEYINPUT55), .B(KEYINPUT83), .Z(n703) );
  XNOR2_X1 U762 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n702) );
  XNOR2_X1 U763 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U764 ( .A(n705), .B(n704), .ZN(n707) );
  XNOR2_X1 U765 ( .A(n709), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U766 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n711) );
  NAND2_X1 U767 ( .A1(n722), .A2(G469), .ZN(n710) );
  BUF_X1 U768 ( .A(n712), .Z(n713) );
  NOR2_X1 U769 ( .A1(n724), .A2(n714), .ZN(G54) );
  NAND2_X1 U770 ( .A1(n722), .A2(G475), .ZN(n717) );
  NAND2_X1 U771 ( .A1(G478), .A2(n722), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n724), .A2(n721), .ZN(G63) );
  XOR2_X1 U774 ( .A(KEYINPUT123), .B(n726), .Z(G66) );
  INV_X1 U775 ( .A(G898), .ZN(n729) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n727) );
  XOR2_X1 U777 ( .A(KEYINPUT61), .B(n727), .Z(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n732) );
  NOR2_X1 U779 ( .A1(G953), .A2(n351), .ZN(n731) );
  NOR2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n739) );
  NOR2_X1 U781 ( .A1(G898), .A2(n733), .ZN(n737) );
  XOR2_X1 U782 ( .A(n735), .B(n734), .Z(n736) );
  NOR2_X1 U783 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U784 ( .A(n739), .B(n738), .Z(G69) );
  XOR2_X1 U785 ( .A(n740), .B(KEYINPUT124), .Z(n741) );
  XNOR2_X1 U786 ( .A(n742), .B(n741), .ZN(n745) );
  NOR2_X1 U787 ( .A1(G953), .A2(n743), .ZN(n744) );
  XNOR2_X1 U788 ( .A(n744), .B(KEYINPUT125), .ZN(n749) );
  XNOR2_X1 U789 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U790 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U791 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U792 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U793 ( .A(n750), .B(G131), .Z(G33) );
  XNOR2_X1 U794 ( .A(G122), .B(KEYINPUT126), .ZN(n751) );
  XNOR2_X1 U795 ( .A(G119), .B(n752), .ZN(G21) );
  XNOR2_X1 U796 ( .A(G134), .B(n753), .ZN(G36) );
  XOR2_X1 U797 ( .A(G137), .B(n754), .Z(G39) );
endmodule

