

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751;

  XOR2_X1 U368 ( .A(G140), .B(G107), .Z(n485) );
  XNOR2_X1 U369 ( .A(G113), .B(G131), .ZN(n451) );
  INV_X1 U370 ( .A(G104), .ZN(n409) );
  NAND2_X2 U371 ( .A1(n352), .A2(n372), .ZN(n346) );
  AND2_X2 U372 ( .A1(n356), .A2(n354), .ZN(n359) );
  XNOR2_X2 U373 ( .A(n346), .B(n544), .ZN(n676) );
  AND2_X2 U374 ( .A1(n376), .A2(n377), .ZN(n362) );
  XNOR2_X2 U375 ( .A(G902), .B(KEYINPUT15), .ZN(n599) );
  OR2_X2 U376 ( .A1(n540), .A2(n512), .ZN(n374) );
  XNOR2_X2 U377 ( .A(n572), .B(n368), .ZN(n434) );
  XNOR2_X1 U378 ( .A(G116), .B(KEYINPUT95), .ZN(n492) );
  XNOR2_X1 U379 ( .A(G122), .B(KEYINPUT98), .ZN(n454) );
  INV_X1 U380 ( .A(G146), .ZN(n414) );
  XNOR2_X1 U381 ( .A(KEYINPUT10), .B(G140), .ZN(n449) );
  BUF_X1 U382 ( .A(G128), .Z(n654) );
  NAND2_X2 U383 ( .A1(n383), .A2(n380), .ZN(n572) );
  AND2_X2 U384 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X2 U385 ( .A1(n513), .A2(n514), .ZN(n515) );
  NAND2_X2 U386 ( .A1(n362), .A2(n374), .ZN(n514) );
  INV_X4 U387 ( .A(G953), .ZN(n741) );
  XNOR2_X1 U388 ( .A(n596), .B(KEYINPUT79), .ZN(n678) );
  NOR2_X1 U389 ( .A1(n543), .A2(n542), .ZN(n373) );
  XNOR2_X1 U390 ( .A(n516), .B(KEYINPUT68), .ZN(n682) );
  OR2_X1 U391 ( .A1(n552), .A2(n553), .ZN(n516) );
  INV_X1 U392 ( .A(G902), .ZN(n505) );
  INV_X1 U393 ( .A(KEYINPUT72), .ZN(n360) );
  BUF_X1 U394 ( .A(n678), .Z(n740) );
  NAND2_X1 U395 ( .A1(n358), .A2(n360), .ZN(n357) );
  OR2_X1 U396 ( .A1(n524), .A2(n525), .ZN(n526) );
  XNOR2_X1 U397 ( .A(n373), .B(KEYINPUT80), .ZN(n372) );
  AND2_X1 U398 ( .A1(n355), .A2(n523), .ZN(n354) );
  AND2_X1 U399 ( .A1(n748), .A2(KEYINPUT44), .ZN(n543) );
  INV_X1 U400 ( .A(n748), .ZN(n402) );
  XNOR2_X1 U401 ( .A(n387), .B(n566), .ZN(n751) );
  NOR2_X1 U402 ( .A1(n577), .A2(n369), .ZN(n669) );
  AND2_X1 U403 ( .A1(n400), .A2(n562), .ZN(n365) );
  XNOR2_X1 U404 ( .A(n399), .B(KEYINPUT92), .ZN(n562) );
  AND2_X1 U405 ( .A1(n563), .A2(n401), .ZN(n400) );
  XOR2_X1 U406 ( .A(KEYINPUT107), .B(n568), .Z(n662) );
  INV_X1 U407 ( .A(n602), .ZN(n349) );
  XOR2_X1 U408 ( .A(KEYINPUT66), .B(n601), .Z(n602) );
  XNOR2_X2 U409 ( .A(G116), .B(G107), .ZN(n420) );
  XNOR2_X1 U410 ( .A(KEYINPUT23), .B(G110), .ZN(n398) );
  XNOR2_X2 U411 ( .A(KEYINPUT99), .B(KEYINPUT11), .ZN(n453) );
  XNOR2_X2 U412 ( .A(KEYINPUT85), .B(G110), .ZN(n410) );
  XNOR2_X2 U413 ( .A(KEYINPUT67), .B(G101), .ZN(n408) );
  XOR2_X2 U414 ( .A(G104), .B(G143), .Z(n452) );
  NOR2_X1 U415 ( .A1(G953), .A2(G237), .ZN(n495) );
  XOR2_X2 U416 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n493) );
  BUF_X2 U417 ( .A(n629), .Z(n638) );
  AND2_X2 U418 ( .A1(n348), .A2(n347), .ZN(n629) );
  INV_X1 U419 ( .A(n674), .ZN(n347) );
  NAND2_X1 U420 ( .A1(n350), .A2(n349), .ZN(n348) );
  INV_X1 U421 ( .A(n603), .ZN(n350) );
  NAND2_X1 U422 ( .A1(n748), .A2(n360), .ZN(n355) );
  XNOR2_X2 U423 ( .A(n404), .B(KEYINPUT35), .ZN(n748) );
  NAND2_X1 U424 ( .A1(n353), .A2(n526), .ZN(n352) );
  NAND2_X1 U425 ( .A1(n359), .A2(n357), .ZN(n353) );
  NAND2_X1 U426 ( .A1(n403), .A2(n361), .ZN(n356) );
  XNOR2_X1 U427 ( .A(n524), .B(KEYINPUT81), .ZN(n403) );
  XNOR2_X2 U428 ( .A(n515), .B(KEYINPUT82), .ZN(n524) );
  XNOR2_X2 U429 ( .A(n498), .B(n728), .ZN(n482) );
  XNOR2_X2 U430 ( .A(n736), .B(n408), .ZN(n498) );
  XNOR2_X2 U431 ( .A(n435), .B(KEYINPUT4), .ZN(n736) );
  XNOR2_X2 U432 ( .A(G143), .B(G128), .ZN(n435) );
  INV_X1 U433 ( .A(n403), .ZN(n358) );
  AND2_X1 U434 ( .A1(n402), .A2(KEYINPUT72), .ZN(n361) );
  NAND2_X1 U435 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U436 ( .A1(n425), .A2(n386), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n398), .B(n654), .ZN(n397) );
  XNOR2_X1 U438 ( .A(n471), .B(n396), .ZN(n395) );
  INV_X1 U439 ( .A(KEYINPUT24), .ZN(n471) );
  INV_X1 U440 ( .A(G119), .ZN(n396) );
  XNOR2_X1 U441 ( .A(n565), .B(KEYINPUT39), .ZN(n595) );
  XNOR2_X1 U442 ( .A(n465), .B(n464), .ZN(n529) );
  XNOR2_X1 U443 ( .A(n463), .B(G475), .ZN(n464) );
  OR2_X1 U444 ( .A1(n511), .A2(n512), .ZN(n378) );
  AND2_X1 U445 ( .A1(n391), .A2(n594), .ZN(n390) );
  NAND2_X1 U446 ( .A1(n585), .A2(KEYINPUT48), .ZN(n391) );
  INV_X1 U447 ( .A(KEYINPUT83), .ZN(n386) );
  NAND2_X1 U448 ( .A1(n425), .A2(n386), .ZN(n384) );
  INV_X1 U449 ( .A(G237), .ZN(n423) );
  XNOR2_X1 U450 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n412) );
  INV_X1 U451 ( .A(KEYINPUT0), .ZN(n370) );
  XNOR2_X1 U452 ( .A(n504), .B(n503), .ZN(n623) );
  NOR2_X1 U453 ( .A1(n682), .A2(n557), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n623), .B(KEYINPUT62), .ZN(n624) );
  XNOR2_X1 U455 ( .A(n473), .B(n394), .ZN(n476) );
  XNOR2_X1 U456 ( .A(n397), .B(n395), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U458 ( .A(n617), .B(n616), .ZN(n618) );
  OR2_X1 U459 ( .A1(n741), .A2(G952), .ZN(n633) );
  NAND2_X1 U460 ( .A1(n595), .A2(n568), .ZN(n387) );
  INV_X1 U461 ( .A(n582), .ZN(n405) );
  AND2_X1 U462 ( .A1(n378), .A2(n553), .ZN(n377) );
  XNOR2_X1 U463 ( .A(n450), .B(n449), .ZN(n474) );
  OR2_X1 U464 ( .A1(n551), .A2(n433), .ZN(n363) );
  NOR2_X1 U465 ( .A1(n585), .A2(KEYINPUT48), .ZN(n364) );
  XNOR2_X1 U466 ( .A(KEYINPUT34), .B(n522), .ZN(n366) );
  NAND2_X1 U467 ( .A1(n424), .A2(G210), .ZN(n367) );
  XOR2_X1 U468 ( .A(KEYINPUT73), .B(KEYINPUT19), .Z(n368) );
  XNOR2_X1 U469 ( .A(n557), .B(KEYINPUT1), .ZN(n369) );
  XNOR2_X1 U470 ( .A(n557), .B(KEYINPUT1), .ZN(n681) );
  XNOR2_X2 U471 ( .A(n371), .B(n370), .ZN(n520) );
  AND2_X2 U472 ( .A1(n434), .A2(n363), .ZN(n371) );
  BUF_X1 U473 ( .A(n435), .Z(n436) );
  NOR2_X2 U474 ( .A1(n520), .A2(n470), .ZN(n407) );
  XNOR2_X2 U475 ( .A(n375), .B(KEYINPUT32), .ZN(n513) );
  NAND2_X1 U476 ( .A1(n540), .A2(n510), .ZN(n375) );
  XNOR2_X2 U477 ( .A(n407), .B(KEYINPUT22), .ZN(n540) );
  NAND2_X1 U478 ( .A1(n540), .A2(n379), .ZN(n376) );
  AND2_X1 U479 ( .A1(n511), .A2(n512), .ZN(n379) );
  INV_X1 U480 ( .A(n545), .ZN(n382) );
  NAND2_X1 U481 ( .A1(n545), .A2(n386), .ZN(n385) );
  INV_X1 U482 ( .A(n434), .ZN(n579) );
  XNOR2_X2 U483 ( .A(n491), .B(n490), .ZN(n557) );
  NAND2_X1 U484 ( .A1(n750), .A2(n751), .ZN(n567) );
  NOR2_X2 U485 ( .A1(n389), .A2(n388), .ZN(n606) );
  AND2_X1 U486 ( .A1(n586), .A2(KEYINPUT48), .ZN(n388) );
  NAND2_X1 U487 ( .A1(n392), .A2(n390), .ZN(n389) );
  NAND2_X1 U488 ( .A1(n393), .A2(n364), .ZN(n392) );
  INV_X1 U489 ( .A(n586), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n606), .A2(n671), .ZN(n596) );
  INV_X1 U491 ( .A(n564), .ZN(n401) );
  NAND2_X1 U492 ( .A1(n366), .A2(n405), .ZN(n404) );
  XNOR2_X2 U493 ( .A(n406), .B(n367), .ZN(n545) );
  NAND2_X1 U494 ( .A1(n614), .A2(n599), .ZN(n406) );
  XNOR2_X1 U495 ( .A(n567), .B(KEYINPUT46), .ZN(n586) );
  INV_X1 U496 ( .A(n672), .ZN(n594) );
  BUF_X1 U497 ( .A(n498), .Z(n499) );
  XNOR2_X1 U498 ( .A(n500), .B(n499), .ZN(n504) );
  NOR2_X1 U499 ( .A1(n571), .A2(n570), .ZN(n587) );
  XNOR2_X1 U500 ( .A(n410), .B(n409), .ZN(n728) );
  NAND2_X1 U501 ( .A1(n741), .A2(G224), .ZN(n411) );
  XNOR2_X1 U502 ( .A(n411), .B(KEYINPUT74), .ZN(n413) );
  XNOR2_X1 U503 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U504 ( .A(n414), .B(G125), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n415), .B(n450), .ZN(n416) );
  XNOR2_X1 U506 ( .A(n482), .B(n416), .ZN(n422) );
  XOR2_X1 U507 ( .A(KEYINPUT3), .B(G119), .Z(n418) );
  XNOR2_X1 U508 ( .A(KEYINPUT71), .B(G113), .ZN(n417) );
  XNOR2_X1 U509 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U510 ( .A(KEYINPUT86), .B(n419), .Z(n502) );
  XNOR2_X1 U511 ( .A(n420), .B(G122), .ZN(n438) );
  XNOR2_X1 U512 ( .A(n438), .B(KEYINPUT16), .ZN(n421) );
  XNOR2_X1 U513 ( .A(n502), .B(n421), .ZN(n730) );
  XNOR2_X1 U514 ( .A(n422), .B(n730), .ZN(n614) );
  NAND2_X1 U515 ( .A1(n505), .A2(n423), .ZN(n424) );
  NAND2_X1 U516 ( .A1(n424), .A2(G214), .ZN(n697) );
  INV_X1 U517 ( .A(n697), .ZN(n425) );
  NAND2_X1 U518 ( .A1(G234), .A2(G237), .ZN(n426) );
  XNOR2_X1 U519 ( .A(n426), .B(KEYINPUT14), .ZN(n428) );
  NAND2_X1 U520 ( .A1(n428), .A2(G952), .ZN(n427) );
  XOR2_X1 U521 ( .A(KEYINPUT87), .B(n427), .Z(n711) );
  NOR2_X1 U522 ( .A1(n711), .A2(G953), .ZN(n551) );
  NAND2_X1 U523 ( .A1(G902), .A2(n428), .ZN(n429) );
  XOR2_X1 U524 ( .A(KEYINPUT88), .B(n429), .Z(n430) );
  NAND2_X1 U525 ( .A1(G953), .A2(n430), .ZN(n548) );
  NOR2_X1 U526 ( .A1(G898), .A2(n548), .ZN(n432) );
  INV_X1 U527 ( .A(KEYINPUT89), .ZN(n431) );
  XNOR2_X1 U528 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U529 ( .A(n436), .B(KEYINPUT7), .ZN(n437) );
  XNOR2_X1 U530 ( .A(n438), .B(n437), .ZN(n445) );
  XOR2_X1 U531 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n440) );
  XNOR2_X1 U532 ( .A(G134), .B(KEYINPUT101), .ZN(n439) );
  XNOR2_X1 U533 ( .A(n440), .B(n439), .ZN(n443) );
  NAND2_X1 U534 ( .A1(G234), .A2(n741), .ZN(n441) );
  XOR2_X1 U535 ( .A(KEYINPUT8), .B(n441), .Z(n472) );
  NAND2_X1 U536 ( .A1(G217), .A2(n472), .ZN(n442) );
  XNOR2_X1 U537 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n635) );
  NOR2_X1 U539 ( .A1(G902), .A2(n635), .ZN(n446) );
  XOR2_X1 U540 ( .A(n446), .B(KEYINPUT103), .Z(n448) );
  INV_X1 U541 ( .A(G478), .ZN(n447) );
  XNOR2_X1 U542 ( .A(n448), .B(n447), .ZN(n528) );
  INV_X1 U543 ( .A(n528), .ZN(n530) );
  XNOR2_X1 U544 ( .A(n452), .B(n451), .ZN(n457) );
  INV_X1 U545 ( .A(n453), .ZN(n455) );
  XNOR2_X1 U546 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U547 ( .A(n457), .B(n456), .Z(n461) );
  XOR2_X1 U548 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n459) );
  NAND2_X1 U549 ( .A1(G214), .A2(n495), .ZN(n458) );
  XNOR2_X1 U550 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U551 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n474), .B(n462), .ZN(n608) );
  NOR2_X1 U553 ( .A1(G902), .A2(n608), .ZN(n465) );
  XNOR2_X1 U554 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n463) );
  INV_X1 U555 ( .A(n529), .ZN(n527) );
  NAND2_X1 U556 ( .A1(n530), .A2(n527), .ZN(n700) );
  NAND2_X1 U557 ( .A1(G234), .A2(n599), .ZN(n466) );
  XNOR2_X1 U558 ( .A(KEYINPUT20), .B(n466), .ZN(n477) );
  NAND2_X1 U559 ( .A1(n477), .A2(G221), .ZN(n469) );
  INV_X1 U560 ( .A(KEYINPUT91), .ZN(n467) );
  XNOR2_X1 U561 ( .A(n467), .B(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U562 ( .A(n469), .B(n468), .ZN(n552) );
  OR2_X1 U563 ( .A1(n700), .A2(n552), .ZN(n470) );
  NAND2_X1 U564 ( .A1(n472), .A2(G221), .ZN(n473) );
  XNOR2_X1 U565 ( .A(G137), .B(n474), .ZN(n475) );
  XNOR2_X1 U566 ( .A(n476), .B(n475), .ZN(n630) );
  NAND2_X1 U567 ( .A1(n630), .A2(n505), .ZN(n481) );
  NAND2_X1 U568 ( .A1(n477), .A2(G217), .ZN(n479) );
  XNOR2_X1 U569 ( .A(KEYINPUT90), .B(KEYINPUT25), .ZN(n478) );
  XNOR2_X1 U570 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U571 ( .A(n481), .B(n480), .ZN(n553) );
  XNOR2_X1 U572 ( .A(n553), .B(KEYINPUT105), .ZN(n684) );
  BUF_X1 U573 ( .A(n482), .Z(n483) );
  NAND2_X1 U574 ( .A1(G227), .A2(n741), .ZN(n484) );
  XNOR2_X1 U575 ( .A(n485), .B(n484), .ZN(n487) );
  XOR2_X2 U576 ( .A(G137), .B(G134), .Z(n486) );
  XNOR2_X1 U577 ( .A(G131), .B(n486), .ZN(n738) );
  XNOR2_X1 U578 ( .A(G146), .B(n738), .ZN(n501) );
  XNOR2_X1 U579 ( .A(n487), .B(n501), .ZN(n488) );
  XNOR2_X1 U580 ( .A(n483), .B(n488), .ZN(n641) );
  OR2_X1 U581 ( .A1(n641), .A2(G902), .ZN(n491) );
  XNOR2_X1 U582 ( .A(G469), .B(KEYINPUT70), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n489), .B(KEYINPUT69), .ZN(n490) );
  NOR2_X1 U584 ( .A1(n684), .A2(n369), .ZN(n509) );
  XNOR2_X1 U585 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U586 ( .A(KEYINPUT93), .B(n494), .Z(n497) );
  NAND2_X1 U587 ( .A1(n495), .A2(G210), .ZN(n496) );
  XNOR2_X1 U588 ( .A(n497), .B(n496), .ZN(n500) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n623), .A2(n505), .ZN(n506) );
  XNOR2_X2 U591 ( .A(n506), .B(G472), .ZN(n688) );
  XNOR2_X1 U592 ( .A(n688), .B(KEYINPUT6), .ZN(n570) );
  INV_X1 U593 ( .A(KEYINPUT75), .ZN(n507) );
  XNOR2_X1 U594 ( .A(n570), .B(n507), .ZN(n508) );
  AND2_X1 U595 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U596 ( .A(n513), .B(G119), .ZN(G21) );
  INV_X1 U597 ( .A(n688), .ZN(n532) );
  AND2_X1 U598 ( .A1(n369), .A2(n532), .ZN(n511) );
  INV_X1 U599 ( .A(KEYINPUT64), .ZN(n512) );
  XNOR2_X1 U600 ( .A(n514), .B(G110), .ZN(G12) );
  NOR2_X1 U601 ( .A1(n682), .A2(n681), .ZN(n535) );
  INV_X1 U602 ( .A(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U603 ( .A(n535), .B(n517), .ZN(n518) );
  NOR2_X1 U604 ( .A1(n518), .A2(n570), .ZN(n519) );
  XNOR2_X1 U605 ( .A(KEYINPUT33), .B(n519), .ZN(n713) );
  BUF_X1 U606 ( .A(n520), .Z(n521) );
  NOR2_X1 U607 ( .A1(n713), .A2(n521), .ZN(n522) );
  NAND2_X1 U608 ( .A1(n528), .A2(n529), .ZN(n582) );
  INV_X1 U609 ( .A(KEYINPUT44), .ZN(n523) );
  NAND2_X1 U610 ( .A1(KEYINPUT72), .A2(KEYINPUT44), .ZN(n525) );
  NOR2_X2 U611 ( .A1(n528), .A2(n527), .ZN(n568) );
  NOR2_X1 U612 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U613 ( .A(KEYINPUT104), .B(n531), .ZN(n664) );
  NOR2_X1 U614 ( .A1(n568), .A2(n664), .ZN(n703) );
  NAND2_X1 U615 ( .A1(n562), .A2(n532), .ZN(n533) );
  NOR2_X1 U616 ( .A1(n521), .A2(n533), .ZN(n534) );
  XNOR2_X1 U617 ( .A(KEYINPUT96), .B(n534), .ZN(n649) );
  NAND2_X1 U618 ( .A1(n535), .A2(n688), .ZN(n692) );
  NOR2_X1 U619 ( .A1(n521), .A2(n692), .ZN(n536) );
  XOR2_X1 U620 ( .A(KEYINPUT31), .B(n536), .Z(n665) );
  NOR2_X1 U621 ( .A1(n649), .A2(n665), .ZN(n537) );
  NOR2_X1 U622 ( .A1(n703), .A2(n537), .ZN(n541) );
  NAND2_X1 U623 ( .A1(n684), .A2(n570), .ZN(n538) );
  INV_X1 U624 ( .A(n369), .ZN(n588) );
  NOR2_X1 U625 ( .A1(n538), .A2(n588), .ZN(n539) );
  AND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n646) );
  OR2_X1 U627 ( .A1(n541), .A2(n646), .ZN(n542) );
  INV_X1 U628 ( .A(KEYINPUT45), .ZN(n544) );
  BUF_X1 U629 ( .A(n545), .Z(n592) );
  XNOR2_X1 U630 ( .A(n592), .B(KEYINPUT38), .ZN(n698) );
  NAND2_X1 U631 ( .A1(n698), .A2(n697), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n546), .B(KEYINPUT112), .ZN(n702) );
  NOR2_X1 U633 ( .A1(n700), .A2(n702), .ZN(n547) );
  XNOR2_X1 U634 ( .A(n547), .B(KEYINPUT41), .ZN(n712) );
  XOR2_X1 U635 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n556) );
  NOR2_X1 U636 ( .A1(G900), .A2(n548), .ZN(n549) );
  XNOR2_X1 U637 ( .A(n549), .B(KEYINPUT108), .ZN(n550) );
  NOR2_X1 U638 ( .A1(n551), .A2(n550), .ZN(n564) );
  INV_X1 U639 ( .A(n552), .ZN(n685) );
  NAND2_X1 U640 ( .A1(n553), .A2(n685), .ZN(n554) );
  NOR2_X1 U641 ( .A1(n564), .A2(n554), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n569), .A2(n688), .ZN(n555) );
  XNOR2_X1 U643 ( .A(n556), .B(n555), .ZN(n559) );
  INV_X1 U644 ( .A(n557), .ZN(n558) );
  NAND2_X1 U645 ( .A1(n559), .A2(n558), .ZN(n578) );
  NOR2_X1 U646 ( .A1(n712), .A2(n578), .ZN(n560) );
  XOR2_X1 U647 ( .A(KEYINPUT42), .B(n560), .Z(n750) );
  XOR2_X1 U648 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n566) );
  NAND2_X1 U649 ( .A1(n688), .A2(n697), .ZN(n561) );
  XOR2_X1 U650 ( .A(KEYINPUT30), .B(n561), .Z(n563) );
  NAND2_X1 U651 ( .A1(n365), .A2(n698), .ZN(n565) );
  XNOR2_X1 U652 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n569), .A2(n662), .ZN(n571) );
  BUF_X1 U654 ( .A(n572), .Z(n573) );
  INV_X1 U655 ( .A(n573), .ZN(n574) );
  NAND2_X1 U656 ( .A1(n587), .A2(n574), .ZN(n575) );
  XOR2_X1 U657 ( .A(n576), .B(n575), .Z(n577) );
  OR2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n655) );
  OR2_X1 U659 ( .A1(n655), .A2(n703), .ZN(n580) );
  XNOR2_X1 U660 ( .A(KEYINPUT47), .B(n580), .ZN(n581) );
  NOR2_X1 U661 ( .A1(n669), .A2(n581), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n592), .A2(n582), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n365), .A2(n583), .ZN(n658) );
  NAND2_X1 U664 ( .A1(n584), .A2(n658), .ZN(n585) );
  XNOR2_X1 U665 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n587), .A2(n697), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U668 ( .A(n591), .B(n590), .Z(n593) );
  NOR2_X1 U669 ( .A1(n593), .A2(n382), .ZN(n672) );
  NAND2_X1 U670 ( .A1(n595), .A2(n664), .ZN(n671) );
  INV_X1 U671 ( .A(n599), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n678), .A2(n597), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n676), .A2(n598), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT78), .B(n599), .Z(n600) );
  NAND2_X1 U675 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  NAND2_X1 U676 ( .A1(KEYINPUT2), .A2(n671), .ZN(n604) );
  XOR2_X1 U677 ( .A(KEYINPUT76), .B(n604), .Z(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n679) );
  NOR2_X1 U679 ( .A1(n676), .A2(n679), .ZN(n674) );
  NAND2_X1 U680 ( .A1(n629), .A2(G475), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n607) );
  XNOR2_X1 U682 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n611), .A2(n633), .ZN(n613) );
  INV_X1 U684 ( .A(KEYINPUT60), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(G60) );
  NAND2_X1 U686 ( .A1(n629), .A2(G210), .ZN(n619) );
  BUF_X1 U687 ( .A(n614), .Z(n617) );
  XNOR2_X1 U688 ( .A(KEYINPUT77), .B(KEYINPUT54), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT55), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n620), .A2(n633), .ZN(n622) );
  INV_X1 U692 ( .A(KEYINPUT56), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(G51) );
  NAND2_X1 U694 ( .A1(n629), .A2(G472), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n626), .A2(n633), .ZN(n628) );
  XNOR2_X1 U697 ( .A(KEYINPUT84), .B(KEYINPUT63), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(G57) );
  NAND2_X1 U699 ( .A1(n638), .A2(G217), .ZN(n632) );
  XOR2_X1 U700 ( .A(KEYINPUT124), .B(n630), .Z(n631) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(n634) );
  INV_X1 U702 ( .A(n633), .ZN(n644) );
  NOR2_X1 U703 ( .A1(n634), .A2(n644), .ZN(G66) );
  NAND2_X1 U704 ( .A1(n638), .A2(G478), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X1 U706 ( .A1(n637), .A2(n644), .ZN(G63) );
  NAND2_X1 U707 ( .A1(n638), .A2(G469), .ZN(n643) );
  XNOR2_X1 U708 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT58), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n643), .B(n642), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n645), .A2(n644), .ZN(G54) );
  XOR2_X1 U713 ( .A(G101), .B(n646), .Z(G3) );
  NAND2_X1 U714 ( .A1(n649), .A2(n662), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  XNOR2_X1 U716 ( .A(G104), .B(n648), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n651) );
  NAND2_X1 U718 ( .A1(n649), .A2(n664), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n653) );
  XOR2_X1 U720 ( .A(G107), .B(KEYINPUT115), .Z(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(G9) );
  XOR2_X1 U722 ( .A(n654), .B(KEYINPUT29), .Z(n657) );
  INV_X1 U723 ( .A(n655), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n659), .A2(n664), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(G30) );
  XNOR2_X1 U726 ( .A(G143), .B(n658), .ZN(G45) );
  NAND2_X1 U727 ( .A1(n659), .A2(n662), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT116), .ZN(n661) );
  XNOR2_X1 U729 ( .A(G146), .B(n661), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n662), .A2(n665), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(G113), .ZN(G15) );
  XOR2_X1 U732 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n667) );
  NAND2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U735 ( .A(G116), .B(n668), .ZN(G18) );
  XNOR2_X1 U736 ( .A(n669), .B(G125), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U738 ( .A(G134), .B(n671), .ZN(G36) );
  XNOR2_X1 U739 ( .A(n672), .B(G140), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(KEYINPUT119), .ZN(G42) );
  INV_X1 U741 ( .A(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n674), .A2(n675), .ZN(n720) );
  BUF_X1 U743 ( .A(n676), .Z(n677) );
  NAND2_X1 U744 ( .A1(n740), .A2(n679), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n677), .A2(n680), .ZN(n718) );
  NAND2_X1 U746 ( .A1(n682), .A2(n369), .ZN(n683) );
  XNOR2_X1 U747 ( .A(KEYINPUT50), .B(n683), .ZN(n690) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(n686), .Z(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U752 ( .A(n691), .B(KEYINPUT120), .ZN(n693) );
  NAND2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n695) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(KEYINPUT121), .Z(n694) );
  XNOR2_X1 U755 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n696), .A2(n712), .ZN(n708) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n701), .B(KEYINPUT122), .ZN(n705) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n706), .A2(n713), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n709), .B(KEYINPUT52), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U767 ( .A1(G953), .A2(n714), .ZN(n715) );
  OR2_X1 U768 ( .A1(n716), .A2(n715), .ZN(n717) );
  OR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U770 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U771 ( .A(KEYINPUT53), .B(n721), .ZN(G75) );
  INV_X1 U772 ( .A(n677), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n722), .A2(n741), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n723) );
  XNOR2_X1 U775 ( .A(KEYINPUT61), .B(n723), .ZN(n724) );
  NAND2_X1 U776 ( .A1(n724), .A2(G898), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n734) );
  XNOR2_X1 U778 ( .A(G101), .B(KEYINPUT125), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U780 ( .A(n730), .B(n729), .ZN(n732) );
  NOR2_X1 U781 ( .A1(n741), .A2(G898), .ZN(n731) );
  NOR2_X1 U782 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U783 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n735), .ZN(G69) );
  BUF_X1 U785 ( .A(n736), .Z(n737) );
  XOR2_X1 U786 ( .A(n737), .B(n738), .Z(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(n474), .ZN(n743) );
  XOR2_X1 U788 ( .A(n743), .B(n740), .Z(n742) );
  NAND2_X1 U789 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U790 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U791 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n747), .A2(n746), .ZN(G72) );
  XNOR2_X1 U794 ( .A(G122), .B(n748), .ZN(n749) );
  XNOR2_X1 U795 ( .A(n749), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U796 ( .A(G137), .B(n750), .ZN(G39) );
  XNOR2_X1 U797 ( .A(n751), .B(G131), .ZN(G33) );
endmodule

