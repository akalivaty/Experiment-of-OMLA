//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n438, new_n439, new_n440, new_n444, new_n445, new_n446, new_n452,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n438));
  OR2_X1    g013(.A1(new_n438), .A2(G69), .ZN(new_n439));
  NAND2_X1  g014(.A1(new_n438), .A2(G69), .ZN(new_n440));
  NAND2_X1  g015(.A1(new_n439), .A2(new_n440), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n444));
  OR2_X1    g019(.A1(new_n444), .A2(G108), .ZN(new_n445));
  NAND2_X1  g020(.A1(new_n444), .A2(G108), .ZN(new_n446));
  NAND2_X1  g021(.A1(new_n445), .A2(new_n446), .ZN(G238));
  NAND4_X1  g022(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g023(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g024(.A(G452), .Z(G391));
  AND2_X1   g025(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g028(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n470), .B1(new_n474), .B2(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n480), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n477), .A2(new_n479), .A3(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n477), .A2(new_n479), .A3(G138), .A4(new_n473), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(G138), .A3(new_n473), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT68), .A2(G114), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT68), .A2(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n502), .B2(G2105), .ZN(new_n503));
  AND4_X1   g078(.A1(G126), .A2(new_n477), .A3(new_n479), .A4(G2105), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT70), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(new_n508), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  AND2_X1   g090(.A1(G75), .A2(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n509), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n512), .B1(new_n508), .B2(G651), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n510), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n518), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(G88), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n518), .A2(G62), .A3(G651), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n511), .A2(new_n513), .ZN(new_n529));
  AND4_X1   g104(.A1(KEYINPUT71), .A2(new_n529), .A3(new_n519), .A4(new_n518), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT71), .B1(new_n514), .B2(new_n518), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n514), .A2(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n533), .A2(new_n534), .A3(new_n536), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND3_X1  g115(.A1(new_n524), .A2(G90), .A3(new_n525), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n510), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND3_X1  g121(.A1(new_n524), .A2(G81), .A3(new_n525), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n514), .A2(G43), .A3(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT72), .ZN(G188));
  NAND2_X1  g134(.A1(new_n532), .A2(G91), .ZN(new_n560));
  INV_X1    g135(.A(new_n518), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  INV_X1    g137(.A(G78), .ZN(new_n563));
  INV_X1    g138(.A(G543), .ZN(new_n564));
  OAI22_X1  g139(.A1(new_n561), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  OAI221_X1 g142(.A(new_n567), .B1(new_n563), .B2(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(G651), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n514), .A2(G53), .A3(G543), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n560), .A2(new_n569), .A3(new_n573), .A4(new_n575), .ZN(G299));
  NAND3_X1  g151(.A1(new_n517), .A2(new_n526), .A3(new_n527), .ZN(G303));
  NAND3_X1  g152(.A1(new_n524), .A2(G87), .A3(new_n525), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n535), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n524), .A2(G86), .A3(new_n525), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n535), .A2(G48), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n510), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(G305));
  NAND3_X1  g161(.A1(new_n524), .A2(G85), .A3(new_n525), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n535), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n510), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n532), .A2(new_n593), .A3(G92), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n524), .A2(new_n525), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT10), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n561), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n535), .A2(G54), .B1(new_n600), .B2(G651), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n594), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n592), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n552), .ZN(G323));
  XOR2_X1   g188(.A(G323), .B(KEYINPUT75), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n485), .A2(G2104), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n485), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n487), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2096), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT76), .Z(G156));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT78), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT79), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AND2_X1   g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n638), .A2(new_n642), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR3_X1    g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(KEYINPUT81), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n652), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n652), .A2(new_n653), .ZN(new_n660));
  MUX2_X1   g235(.A(new_n660), .B(new_n652), .S(new_n654), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n656), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n619), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n668), .A2(new_n671), .A3(new_n673), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n676), .B(new_n677), .C1(new_n675), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT82), .B(G1986), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR3_X1    g262(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n684), .B2(new_n685), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  AND2_X1   g265(.A1(KEYINPUT83), .A2(G16), .ZN(new_n691));
  NOR2_X1   g266(.A1(KEYINPUT83), .A2(G16), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G20), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT100), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT23), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G299), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1956), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n473), .ZN(new_n699));
  INV_X1    g274(.A(G139), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n699), .A2(KEYINPUT88), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT88), .B1(new_n699), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(G115), .A2(G2104), .ZN(new_n703));
  INV_X1    g278(.A(G127), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n480), .B2(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n701), .A2(new_n702), .B1(G2105), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT25), .Z(new_n708));
  NAND3_X1  g283(.A1(new_n706), .A2(KEYINPUT89), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(KEYINPUT89), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G29), .B2(G33), .ZN(new_n714));
  INV_X1    g289(.A(G2072), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n698), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT96), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G5), .B2(G16), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n717), .A2(G5), .A3(G16), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(G301), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G16), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G286), .B2(new_n720), .ZN(new_n725));
  INV_X1    g300(.A(G1966), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT95), .Z(new_n728));
  NOR3_X1   g303(.A1(new_n716), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(G160), .A2(G29), .B1(KEYINPUT91), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(KEYINPUT91), .B2(new_n733), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(G2084), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(G2084), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT98), .B(G2078), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G27), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G164), .B2(new_n739), .ZN(new_n741));
  MUX2_X1   g316(.A(new_n740), .B(new_n741), .S(KEYINPUT97), .Z(new_n742));
  AOI22_X1  g317(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n739), .A2(G26), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n485), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n487), .A2(G128), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n739), .ZN(new_n751));
  MUX2_X1   g326(.A(new_n744), .B(new_n751), .S(KEYINPUT28), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT87), .B(G2067), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT30), .B(G28), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n755), .A2(new_n739), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n625), .B2(new_n739), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  OR2_X1    g335(.A1(new_n742), .A2(new_n738), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n743), .A2(new_n754), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n720), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n602), .B2(new_n720), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT86), .ZN(new_n765));
  INV_X1    g340(.A(G1348), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n739), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n487), .A2(G129), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT26), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n467), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n771), .B(new_n773), .C1(new_n774), .C2(G2105), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT92), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT92), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n770), .B1(new_n779), .B2(new_n739), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT93), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT27), .B(G1996), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n693), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n552), .B2(new_n693), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n729), .A2(new_n769), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n725), .A2(new_n726), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n714), .A2(new_n715), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n739), .A2(G35), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G162), .B2(new_n739), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT99), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT29), .B(G2090), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n796), .B(new_n797), .Z(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n790), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT85), .B(KEYINPUT36), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n485), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n487), .A2(G119), .ZN(new_n804));
  NOR2_X1   g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(G29), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT84), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G23), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n578), .A2(new_n580), .A3(new_n579), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT33), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1976), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n693), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n693), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n814), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n814), .A2(new_n819), .A3(KEYINPUT34), .A4(new_n823), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n810), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G290), .B(G24), .S(new_n693), .Z(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n802), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n831), .A3(new_n802), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n800), .B1(new_n833), .B2(new_n834), .ZN(G311));
  NOR4_X1   g410(.A1(new_n787), .A2(new_n792), .A3(new_n798), .A4(new_n789), .ZN(new_n836));
  INV_X1    g411(.A(new_n834), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n832), .ZN(G150));
  NAND3_X1  g413(.A1(new_n524), .A2(G93), .A3(new_n525), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n510), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n535), .A2(G55), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n552), .A2(new_n843), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n847), .A2(new_n841), .A3(new_n839), .A4(new_n842), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n602), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n845), .B1(new_n853), .B2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT101), .Z(G145));
  INV_X1    g430(.A(G142), .ZN(new_n856));
  NOR2_X1   g431(.A1(G106), .A2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n699), .A2(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G130), .B2(new_n487), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n617), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n807), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT102), .B1(new_n503), .B2(new_n504), .ZN(new_n864));
  OR2_X1    g439(.A1(KEYINPUT68), .A2(G114), .ZN(new_n865));
  NAND2_X1  g440(.A1(KEYINPUT68), .A2(G114), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(G2105), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n499), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n749), .B(KEYINPUT103), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n778), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n778), .A2(new_n874), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n498), .B(new_n873), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT104), .B1(new_n710), .B2(new_n711), .ZN(new_n878));
  INV_X1    g453(.A(new_n711), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n709), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n778), .A2(new_n874), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n871), .B1(new_n869), .B2(new_n870), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n498), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n778), .A2(new_n874), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n877), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n877), .A2(new_n888), .B1(new_n880), .B2(new_n712), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n863), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G162), .B(G160), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n625), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n888), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n886), .B1(new_n883), .B2(new_n887), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n881), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n889), .A3(new_n862), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n890), .A2(new_n891), .A3(new_n863), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n862), .B1(new_n898), .B2(new_n889), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT105), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n907), .B(new_n894), .C1(new_n903), .C2(new_n904), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n843), .A2(new_n605), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n587), .A2(new_n588), .ZN(new_n913));
  AOI21_X1  g488(.A(G288), .B1(new_n913), .B2(new_n590), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n816), .A2(G290), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G166), .B(G305), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(G288), .A3(new_n590), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n816), .A2(G290), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G303), .B(G305), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n922), .B(new_n912), .C1(new_n914), .C2(new_n915), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(KEYINPUT108), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n926), .B(new_n927), .Z(new_n928));
  NAND3_X1  g503(.A1(new_n594), .A2(new_n597), .A3(new_n601), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(G299), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(KEYINPUT106), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  INV_X1    g512(.A(new_n931), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n929), .A2(G299), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(KEYINPUT41), .A3(new_n931), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n611), .B(new_n849), .ZN(new_n943));
  MUX2_X1   g518(.A(new_n936), .B(new_n942), .S(new_n943), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n928), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n911), .B1(new_n945), .B2(new_n605), .ZN(G295));
  OAI21_X1  g521(.A(new_n911), .B1(new_n945), .B2(new_n605), .ZN(G331));
  NAND2_X1  g522(.A1(G171), .A2(KEYINPUT109), .ZN(new_n948));
  NAND2_X1  g523(.A1(G168), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(G301), .A2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n846), .A2(new_n848), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n951), .B1(new_n846), .B2(new_n848), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n951), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n839), .A2(new_n842), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n847), .B1(new_n956), .B2(new_n841), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n550), .B1(new_n532), .B2(G81), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n843), .B1(new_n958), .B2(new_n549), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G286), .B1(KEYINPUT109), .B2(G171), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n846), .A2(new_n848), .A3(new_n951), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n940), .A2(new_n954), .A3(new_n941), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n932), .B1(new_n954), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n924), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(KEYINPUT110), .A3(new_n901), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n921), .A2(new_n923), .ZN(new_n969));
  INV_X1    g544(.A(new_n932), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n952), .A2(new_n953), .A3(new_n949), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n954), .A2(new_n963), .A3(new_n940), .A4(new_n941), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n975), .B2(G37), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n973), .A2(new_n969), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n967), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n936), .B1(new_n963), .B2(new_n954), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n924), .B1(new_n981), .B2(new_n964), .ZN(new_n982));
  AND4_X1   g557(.A1(KEYINPUT43), .A2(new_n982), .A3(new_n901), .A4(new_n977), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT44), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n982), .A2(new_n979), .A3(new_n901), .A4(new_n977), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n984), .A2(new_n989), .ZN(G397));
  AOI21_X1  g565(.A(G1384), .B1(new_n873), .B2(new_n498), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  AOI211_X1 g569(.A(new_n994), .B(new_n470), .C1(new_n474), .C2(new_n483), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(G1996), .A3(new_n778), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n997), .A2(KEYINPUT112), .A3(G1996), .A4(new_n778), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G2067), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n749), .B(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n778), .B2(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n997), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n807), .B(new_n809), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n997), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n913), .A2(new_n830), .A3(new_n590), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n996), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n582), .A2(new_n583), .A3(new_n682), .A4(new_n585), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1015), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1022));
  INV_X1    g597(.A(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n991), .B2(new_n995), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1017), .A2(KEYINPUT116), .A3(new_n1018), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n816), .A2(G1976), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  NAND2_X1  g604(.A1(G288), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(KEYINPUT115), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1026), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1384), .B1(new_n498), .B2(new_n505), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n995), .B1(KEYINPUT45), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n886), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(new_n993), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n991), .A2(KEYINPUT114), .A3(KEYINPUT45), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n886), .A2(new_n1044), .A3(new_n1039), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n506), .A2(new_n1039), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(new_n995), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1043), .A2(G1971), .B1(G2090), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1050), .B(KEYINPUT55), .Z(new_n1051));
  AND3_X1   g626(.A1(new_n1049), .A2(G8), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1051), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1044), .B1(new_n886), .B2(new_n1039), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n474), .A2(new_n483), .ZN(new_n1055));
  INV_X1    g630(.A(new_n470), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(G40), .A3(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT50), .B(G1384), .C1(new_n498), .C2(new_n505), .ZN(new_n1058));
  NOR4_X1   g633(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .A4(G2090), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(new_n993), .B2(new_n1046), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT114), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1061));
  AND4_X1   g636(.A1(KEYINPUT114), .A2(new_n886), .A3(KEYINPUT45), .A4(new_n1039), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1063), .B2(new_n822), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1053), .B1(new_n1064), .B2(new_n1023), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1068));
  INV_X1    g643(.A(G2090), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(new_n995), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1043), .B2(G1971), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G8), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .A3(new_n1053), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1035), .B(new_n1052), .C1(new_n1067), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n995), .B(new_n1075), .C1(new_n991), .C2(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n726), .ZN(new_n1077));
  INV_X1    g652(.A(G2084), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1045), .A2(new_n1047), .A3(new_n1078), .A4(new_n995), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(G168), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g659(.A(G286), .B1(new_n1084), .B2(KEYINPUT123), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT123), .B1(new_n1080), .B2(G8), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1088), .B2(KEYINPUT122), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1091));
  INV_X1    g666(.A(G2078), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1043), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n722), .B2(new_n1048), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(KEYINPUT53), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1076), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1087), .A2(new_n1099), .A3(new_n1089), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1074), .A2(new_n1091), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1052), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT117), .B1(new_n1072), .B2(new_n1053), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1066), .B(new_n1051), .C1(new_n1071), .C2(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1023), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1107), .A2(KEYINPUT118), .A3(G168), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT118), .B1(new_n1107), .B2(G168), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1102), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1026), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1049), .A2(G8), .ZN(new_n1114));
  OAI221_X1 g689(.A(new_n1112), .B1(new_n1108), .B2(new_n1109), .C1(new_n1051), .C2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1026), .A2(new_n1029), .A3(new_n816), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1016), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(KEYINPUT63), .B1(new_n1024), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1101), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT56), .B(G2072), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1060), .B(new_n1120), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1058), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n995), .B(new_n1122), .C1(new_n991), .C2(new_n1044), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G299), .B(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1040), .A2(new_n1057), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1048), .A2(new_n766), .B1(new_n1131), .B2(new_n1003), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n929), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1048), .A2(new_n766), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1003), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n602), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1130), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(KEYINPUT120), .A3(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI211_X1 g720(.A(G1996), .B(new_n1037), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1040), .B2(new_n1057), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT121), .B(new_n1147), .C1(new_n1040), .C2(new_n1057), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n552), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1132), .A2(new_n929), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1134), .A2(new_n929), .A3(new_n1135), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT60), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI211_X1 g733(.A(KEYINPUT59), .B(new_n552), .C1(new_n1146), .C2(new_n1152), .ZN(new_n1159));
  OR3_X1    g734(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n929), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1140), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1128), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1140), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1161), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1145), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(G301), .B(KEYINPUT54), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1052), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n472), .A2(new_n473), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1175), .B(new_n1096), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n992), .A2(new_n993), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1176), .A2(G40), .A3(new_n1056), .A4(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1095), .A2(new_n1171), .A3(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1173), .A2(new_n1112), .A3(new_n1174), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1169), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1014), .B1(new_n1119), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n807), .A2(new_n809), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1000), .A2(new_n1001), .A3(new_n1006), .A4(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n750), .A2(new_n1003), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n997), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n996), .A2(G1996), .ZN(new_n1188));
  AND2_X1   g763(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1189));
  INV_X1    g764(.A(G1996), .ZN(new_n1190));
  NOR2_X1   g765(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n779), .A2(new_n1004), .A3(new_n1192), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1188), .A2(new_n1189), .B1(new_n996), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT47), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n996), .A2(new_n1011), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT48), .Z(new_n1197));
  NAND4_X1  g772(.A1(new_n1002), .A2(new_n1197), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1187), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1187), .A2(KEYINPUT125), .A3(new_n1195), .A4(new_n1198), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1182), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(new_n986), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1206), .B1(KEYINPUT43), .B2(new_n978), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n465), .B1(new_n688), .B2(new_n689), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n1208), .A2(KEYINPUT126), .A3(new_n649), .A4(new_n665), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n909), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G401), .A2(G227), .ZN(new_n1211));
  AOI21_X1  g785(.A(KEYINPUT126), .B1(new_n1211), .B2(new_n1208), .ZN(new_n1212));
  NOR3_X1   g786(.A1(new_n1207), .A2(new_n1210), .A3(new_n1212), .ZN(G308));
  AND2_X1   g787(.A1(new_n909), .A2(new_n1209), .ZN(new_n1214));
  AND2_X1   g788(.A1(new_n1211), .A2(new_n1208), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n1214), .B(new_n987), .C1(KEYINPUT126), .C2(new_n1215), .ZN(G225));
endmodule


