

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747;

  AND2_X1 U368 ( .A1(n370), .A2(n365), .ZN(n353) );
  AND2_X1 U369 ( .A1(n550), .A2(n549), .ZN(n569) );
  AND2_X1 U370 ( .A1(n567), .A2(n566), .ZN(n568) );
  OR2_X1 U371 ( .A1(n553), .A2(n548), .ZN(n549) );
  AND2_X1 U372 ( .A1(n500), .A2(n499), .ZN(n542) );
  XNOR2_X1 U373 ( .A(n525), .B(n524), .ZN(n543) );
  INV_X1 U374 ( .A(n532), .ZN(n554) );
  INV_X1 U375 ( .A(KEYINPUT0), .ZN(n348) );
  XNOR2_X1 U376 ( .A(n414), .B(n413), .ZN(n456) );
  BUF_X1 U377 ( .A(G110), .Z(n347) );
  NAND2_X1 U378 ( .A1(n532), .A2(n492), .ZN(n495) );
  XNOR2_X2 U379 ( .A(n491), .B(n348), .ZN(n532) );
  INV_X1 U380 ( .A(G953), .ZN(n735) );
  OR2_X2 U381 ( .A1(n746), .A2(KEYINPUT44), .ZN(n551) );
  XNOR2_X2 U382 ( .A(n539), .B(KEYINPUT35), .ZN(n746) );
  NAND2_X2 U383 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U384 ( .A1(n537), .A2(n506), .ZN(n659) );
  AND2_X1 U385 ( .A1(n561), .A2(n659), .ZN(n672) );
  XNOR2_X1 U386 ( .A(KEYINPUT88), .B(G110), .ZN(n358) );
  INV_X1 U387 ( .A(G143), .ZN(n362) );
  OR2_X1 U388 ( .A1(n546), .A2(n541), .ZN(n550) );
  NAND2_X1 U389 ( .A1(n597), .A2(n490), .ZN(n491) );
  OR2_X1 U390 ( .A1(n537), .A2(n506), .ZN(n662) );
  OR2_X1 U391 ( .A1(n642), .A2(G902), .ZN(n422) );
  XNOR2_X1 U392 ( .A(n731), .B(n404), .ZN(n709) );
  XNOR2_X1 U393 ( .A(n415), .B(KEYINPUT95), .ZN(n731) );
  XNOR2_X1 U394 ( .A(n467), .B(n360), .ZN(n415) );
  XNOR2_X1 U395 ( .A(n451), .B(n398), .ZN(n467) );
  XNOR2_X1 U396 ( .A(n362), .B(G128), .ZN(n451) );
  XNOR2_X1 U397 ( .A(n359), .B(n358), .ZN(n455) );
  XNOR2_X1 U398 ( .A(G107), .B(G104), .ZN(n359) );
  XNOR2_X2 U399 ( .A(n587), .B(n484), .ZN(n597) );
  NAND2_X2 U400 ( .A1(n719), .A2(n734), .ZN(n373) );
  XNOR2_X2 U401 ( .A(n571), .B(n570), .ZN(n719) );
  XNOR2_X2 U402 ( .A(n578), .B(n497), .ZN(n530) );
  INV_X1 U403 ( .A(KEYINPUT65), .ZN(n369) );
  NAND2_X1 U404 ( .A1(n371), .A2(n367), .ZN(n366) );
  NAND2_X1 U405 ( .A1(n369), .A2(KEYINPUT2), .ZN(n367) );
  XNOR2_X1 U406 ( .A(n397), .B(n361), .ZN(n360) );
  XNOR2_X1 U407 ( .A(G137), .B(G131), .ZN(n397) );
  XNOR2_X1 U408 ( .A(KEYINPUT4), .B(KEYINPUT71), .ZN(n361) );
  XOR2_X1 U409 ( .A(n347), .B(G119), .Z(n384) );
  XNOR2_X1 U410 ( .A(G128), .B(G137), .ZN(n383) );
  XNOR2_X1 U411 ( .A(G113), .B(G104), .ZN(n428) );
  XNOR2_X1 U412 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U413 ( .A(G143), .B(G131), .ZN(n433) );
  INV_X1 U414 ( .A(KEYINPUT11), .ZN(n435) );
  XNOR2_X1 U415 ( .A(n445), .B(G140), .ZN(n377) );
  XNOR2_X1 U416 ( .A(n441), .B(n440), .ZN(n537) );
  NOR2_X1 U417 ( .A1(n672), .A2(n594), .ZN(n595) );
  INV_X1 U418 ( .A(G237), .ZN(n423) );
  NAND2_X1 U419 ( .A1(n368), .A2(n366), .ZN(n365) );
  NAND2_X1 U420 ( .A1(n373), .A2(n354), .ZN(n370) );
  NAND2_X1 U421 ( .A1(n619), .A2(n369), .ZN(n368) );
  XNOR2_X1 U422 ( .A(KEYINPUT91), .B(KEYINPUT79), .ZN(n448) );
  XNOR2_X1 U423 ( .A(KEYINPUT4), .B(KEYINPUT90), .ZN(n449) );
  XOR2_X1 U424 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n443) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n406) );
  XNOR2_X1 U426 ( .A(n356), .B(KEYINPUT33), .ZN(n533) );
  AND2_X1 U427 ( .A1(n678), .A2(n531), .ZN(n357) );
  XNOR2_X1 U428 ( .A(G116), .B(G107), .ZN(n468) );
  OR2_X1 U429 ( .A1(G902), .A2(n715), .ZN(n475) );
  BUF_X1 U430 ( .A(n501), .Z(n682) );
  XNOR2_X1 U431 ( .A(n388), .B(n387), .ZN(n628) );
  XNOR2_X1 U432 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U433 ( .A(n732), .B(n380), .ZN(n388) );
  XNOR2_X1 U434 ( .A(n438), .B(n437), .ZN(n622) );
  XNOR2_X1 U435 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U436 ( .A(n430), .B(n374), .ZN(n431) );
  XNOR2_X1 U437 ( .A(n403), .B(n402), .ZN(n404) );
  AND2_X1 U438 ( .A1(n625), .A2(G953), .ZN(n718) );
  OR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n349) );
  AND2_X1 U440 ( .A1(n537), .A2(n536), .ZN(n350) );
  XOR2_X1 U441 ( .A(n426), .B(n425), .Z(n351) );
  XOR2_X1 U442 ( .A(n600), .B(KEYINPUT75), .Z(n352) );
  AND2_X1 U443 ( .A1(KEYINPUT65), .A2(n372), .ZN(n354) );
  INV_X1 U444 ( .A(KEYINPUT2), .ZN(n372) );
  AND2_X1 U445 ( .A1(n371), .A2(n369), .ZN(n355) );
  INV_X1 U446 ( .A(n533), .ZN(n675) );
  NAND2_X1 U447 ( .A1(n357), .A2(n530), .ZN(n356) );
  NAND2_X1 U448 ( .A1(n353), .A2(n363), .ZN(n621) );
  NAND2_X1 U449 ( .A1(n364), .A2(n355), .ZN(n363) );
  INV_X1 U450 ( .A(n373), .ZN(n364) );
  INV_X1 U451 ( .A(n373), .ZN(n665) );
  INV_X1 U452 ( .A(n619), .ZN(n371) );
  BUF_X1 U453 ( .A(n483), .Z(n512) );
  XNOR2_X2 U454 ( .A(n457), .B(n456), .ZN(n726) );
  XNOR2_X1 U455 ( .A(KEYINPUT102), .B(KEYINPUT12), .ZN(n374) );
  AND2_X1 U456 ( .A1(n559), .A2(n504), .ZN(n375) );
  INV_X1 U457 ( .A(KEYINPUT85), .ZN(n544) );
  INV_X1 U458 ( .A(n747), .ZN(n582) );
  INV_X1 U459 ( .A(KEYINPUT10), .ZN(n376) );
  OR2_X1 U460 ( .A1(n537), .A2(n536), .ZN(n670) );
  INV_X1 U461 ( .A(KEYINPUT34), .ZN(n534) );
  XNOR2_X1 U462 ( .A(n466), .B(n465), .ZN(n483) );
  XNOR2_X2 U463 ( .A(n399), .B(G125), .ZN(n445) );
  XNOR2_X2 U464 ( .A(n377), .B(n376), .ZN(n732) );
  XOR2_X1 U465 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n379) );
  XNOR2_X1 U466 ( .A(KEYINPUT23), .B(KEYINPUT98), .ZN(n378) );
  XNOR2_X1 U467 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U468 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n382) );
  NAND2_X1 U469 ( .A1(G234), .A2(n735), .ZN(n381) );
  XNOR2_X1 U470 ( .A(n382), .B(n381), .ZN(n472) );
  NAND2_X1 U471 ( .A1(G221), .A2(n472), .ZN(n386) );
  XNOR2_X1 U472 ( .A(n384), .B(n383), .ZN(n385) );
  INV_X1 U473 ( .A(G902), .ZN(n439) );
  NAND2_X1 U474 ( .A1(n628), .A2(n439), .ZN(n393) );
  XOR2_X1 U475 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n390) );
  XNOR2_X1 U476 ( .A(G902), .B(KEYINPUT15), .ZN(n619) );
  NAND2_X1 U477 ( .A1(G234), .A2(n619), .ZN(n389) );
  XNOR2_X1 U478 ( .A(n390), .B(n389), .ZN(n394) );
  NAND2_X1 U479 ( .A1(n394), .A2(G217), .ZN(n391) );
  XNOR2_X1 U480 ( .A(n391), .B(KEYINPUT25), .ZN(n392) );
  XNOR2_X2 U481 ( .A(n393), .B(n392), .ZN(n496) );
  NAND2_X1 U482 ( .A1(n394), .A2(G221), .ZN(n396) );
  XNOR2_X1 U483 ( .A(KEYINPUT100), .B(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U484 ( .A(n396), .B(n395), .ZN(n680) );
  OR2_X2 U485 ( .A1(n496), .A2(n680), .ZN(n555) );
  INV_X1 U486 ( .A(G134), .ZN(n398) );
  XNOR2_X1 U487 ( .A(KEYINPUT69), .B(G101), .ZN(n444) );
  INV_X2 U488 ( .A(G146), .ZN(n399) );
  XNOR2_X1 U489 ( .A(n444), .B(G146), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n455), .B(n419), .ZN(n403) );
  XOR2_X1 U491 ( .A(KEYINPUT96), .B(G140), .Z(n401) );
  NAND2_X1 U492 ( .A1(G227), .A2(n735), .ZN(n400) );
  XNOR2_X1 U493 ( .A(n401), .B(n400), .ZN(n402) );
  NAND2_X1 U494 ( .A1(n709), .A2(n439), .ZN(n405) );
  INV_X1 U495 ( .A(G469), .ZN(n705) );
  XNOR2_X2 U496 ( .A(n405), .B(n705), .ZN(n578) );
  NOR2_X2 U497 ( .A1(n555), .A2(n578), .ZN(n559) );
  XNOR2_X1 U498 ( .A(KEYINPUT14), .B(n406), .ZN(n408) );
  NAND2_X1 U499 ( .A1(G952), .A2(n408), .ZN(n697) );
  NOR2_X1 U500 ( .A1(n697), .A2(G953), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n407), .B(KEYINPUT93), .ZN(n489) );
  NAND2_X1 U502 ( .A1(G902), .A2(n408), .ZN(n485) );
  NOR2_X1 U503 ( .A1(G900), .A2(n485), .ZN(n409) );
  NAND2_X1 U504 ( .A1(n409), .A2(G953), .ZN(n410) );
  NAND2_X1 U505 ( .A1(n489), .A2(n410), .ZN(n504) );
  XNOR2_X1 U506 ( .A(G119), .B(G116), .ZN(n412) );
  XNOR2_X1 U507 ( .A(G113), .B(KEYINPUT72), .ZN(n411) );
  XNOR2_X1 U508 ( .A(n412), .B(n411), .ZN(n414) );
  XNOR2_X1 U509 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U510 ( .A(n415), .B(n456), .ZN(n421) );
  XNOR2_X1 U511 ( .A(KEYINPUT77), .B(n349), .ZN(n432) );
  NAND2_X1 U512 ( .A1(n432), .A2(G210), .ZN(n417) );
  XNOR2_X1 U513 ( .A(KEYINPUT101), .B(KEYINPUT5), .ZN(n416) );
  XNOR2_X1 U514 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U516 ( .A(n421), .B(n420), .ZN(n642) );
  INV_X1 U517 ( .A(G472), .ZN(n640) );
  XNOR2_X2 U518 ( .A(n422), .B(n640), .ZN(n501) );
  NAND2_X1 U519 ( .A1(n439), .A2(n423), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n463), .A2(G214), .ZN(n667) );
  INV_X1 U521 ( .A(n667), .ZN(n482) );
  NOR2_X1 U522 ( .A1(n501), .A2(n482), .ZN(n426) );
  XNOR2_X1 U523 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n424) );
  XNOR2_X1 U524 ( .A(n424), .B(KEYINPUT107), .ZN(n425) );
  NAND2_X1 U525 ( .A1(n375), .A2(n351), .ZN(n427) );
  XNOR2_X1 U526 ( .A(n427), .B(KEYINPUT78), .ZN(n479) );
  XOR2_X1 U527 ( .A(KEYINPUT103), .B(G122), .Z(n429) );
  XNOR2_X1 U528 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U529 ( .A(n732), .B(n431), .ZN(n438) );
  AND2_X1 U530 ( .A1(n432), .A2(G214), .ZN(n434) );
  NAND2_X1 U531 ( .A1(n622), .A2(n439), .ZN(n441) );
  XOR2_X1 U532 ( .A(KEYINPUT13), .B(G475), .Z(n440) );
  NAND2_X1 U533 ( .A1(G224), .A2(n735), .ZN(n442) );
  XNOR2_X1 U534 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U535 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U536 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U537 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U538 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U539 ( .A(n453), .B(n452), .ZN(n458) );
  XNOR2_X1 U540 ( .A(KEYINPUT16), .B(G122), .ZN(n454) );
  XNOR2_X1 U541 ( .A(n455), .B(n454), .ZN(n457) );
  NAND2_X1 U542 ( .A1(n458), .A2(n726), .ZN(n462) );
  INV_X1 U543 ( .A(n458), .ZN(n460) );
  INV_X1 U544 ( .A(n726), .ZN(n459) );
  NAND2_X1 U545 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U546 ( .A1(n462), .A2(n461), .ZN(n633) );
  NAND2_X1 U547 ( .A1(n633), .A2(n619), .ZN(n466) );
  NAND2_X1 U548 ( .A1(n463), .A2(G210), .ZN(n464) );
  XNOR2_X1 U549 ( .A(n464), .B(KEYINPUT92), .ZN(n465) );
  XNOR2_X1 U550 ( .A(n467), .B(G122), .ZN(n471) );
  XNOR2_X1 U551 ( .A(n468), .B(KEYINPUT9), .ZN(n469) );
  XOR2_X1 U552 ( .A(n469), .B(KEYINPUT7), .Z(n470) );
  XNOR2_X1 U553 ( .A(n471), .B(n470), .ZN(n474) );
  NAND2_X1 U554 ( .A1(G217), .A2(n472), .ZN(n473) );
  XOR2_X1 U555 ( .A(n474), .B(n473), .Z(n715) );
  XNOR2_X1 U556 ( .A(G478), .B(n475), .ZN(n536) );
  INV_X1 U557 ( .A(n536), .ZN(n506) );
  NOR2_X1 U558 ( .A1(n512), .A2(n506), .ZN(n476) );
  NAND2_X1 U559 ( .A1(n537), .A2(n476), .ZN(n477) );
  OR2_X1 U560 ( .A1(n479), .A2(n477), .ZN(n602) );
  XNOR2_X1 U561 ( .A(n602), .B(G143), .ZN(G45) );
  INV_X1 U562 ( .A(KEYINPUT38), .ZN(n478) );
  XNOR2_X1 U563 ( .A(n512), .B(n478), .ZN(n573) );
  OR2_X2 U564 ( .A1(n479), .A2(n573), .ZN(n480) );
  XNOR2_X2 U565 ( .A(n480), .B(KEYINPUT39), .ZN(n526) );
  XNOR2_X1 U566 ( .A(n662), .B(KEYINPUT104), .ZN(n561) );
  INV_X1 U567 ( .A(n561), .ZN(n481) );
  NAND2_X1 U568 ( .A1(n526), .A2(n481), .ZN(n615) );
  XNOR2_X1 U569 ( .A(n615), .B(G134), .ZN(G36) );
  OR2_X2 U570 ( .A1(n483), .A2(n482), .ZN(n587) );
  XNOR2_X1 U571 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n484) );
  INV_X1 U572 ( .A(n485), .ZN(n486) );
  NOR2_X1 U573 ( .A1(G898), .A2(n735), .ZN(n727) );
  NAND2_X1 U574 ( .A1(n486), .A2(n727), .ZN(n487) );
  XNOR2_X1 U575 ( .A(n487), .B(KEYINPUT94), .ZN(n488) );
  NAND2_X1 U576 ( .A1(n489), .A2(n488), .ZN(n490) );
  NOR2_X1 U577 ( .A1(n670), .A2(n680), .ZN(n492) );
  XNOR2_X1 U578 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n493), .B(KEYINPUT73), .ZN(n494) );
  XNOR2_X2 U580 ( .A(n495), .B(n494), .ZN(n523) );
  AND2_X1 U581 ( .A1(n523), .A2(n496), .ZN(n500) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n497) );
  INV_X1 U583 ( .A(n530), .ZN(n509) );
  INV_X1 U584 ( .A(n682), .ZN(n498) );
  NOR2_X1 U585 ( .A1(n530), .A2(n498), .ZN(n499) );
  XOR2_X1 U586 ( .A(n347), .B(n542), .Z(G12) );
  XNOR2_X1 U587 ( .A(n501), .B(KEYINPUT6), .ZN(n531) );
  INV_X1 U588 ( .A(n496), .ZN(n502) );
  NOR2_X1 U589 ( .A1(n680), .A2(n502), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n504), .A2(n503), .ZN(n575) );
  INV_X1 U591 ( .A(n575), .ZN(n505) );
  NAND2_X1 U592 ( .A1(n531), .A2(n505), .ZN(n507) );
  NOR2_X1 U593 ( .A1(n507), .A2(n659), .ZN(n586) );
  NAND2_X1 U594 ( .A1(n586), .A2(n667), .ZN(n508) );
  XOR2_X1 U595 ( .A(KEYINPUT106), .B(n508), .Z(n510) );
  NAND2_X1 U596 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U597 ( .A(n511), .B(KEYINPUT43), .ZN(n513) );
  NAND2_X1 U598 ( .A1(n513), .A2(n512), .ZN(n616) );
  XNOR2_X1 U599 ( .A(n616), .B(G140), .ZN(G42) );
  OR2_X1 U600 ( .A1(n530), .A2(n496), .ZN(n514) );
  NOR2_X1 U601 ( .A1(n514), .A2(n531), .ZN(n515) );
  NAND2_X1 U602 ( .A1(n523), .A2(n515), .ZN(n517) );
  INV_X1 U603 ( .A(KEYINPUT105), .ZN(n516) );
  XNOR2_X1 U604 ( .A(n517), .B(n516), .ZN(n565) );
  XNOR2_X1 U605 ( .A(G101), .B(KEYINPUT112), .ZN(n518) );
  XNOR2_X1 U606 ( .A(n565), .B(n518), .ZN(G3) );
  INV_X1 U607 ( .A(n531), .ZN(n519) );
  XNOR2_X1 U608 ( .A(n519), .B(KEYINPUT80), .ZN(n520) );
  AND2_X1 U609 ( .A1(n520), .A2(n530), .ZN(n521) );
  AND2_X1 U610 ( .A1(n496), .A2(n521), .ZN(n522) );
  NAND2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n525) );
  INV_X1 U612 ( .A(KEYINPUT32), .ZN(n524) );
  XOR2_X1 U613 ( .A(n543), .B(G119), .Z(G21) );
  INV_X1 U614 ( .A(n659), .ZN(n657) );
  NAND2_X2 U615 ( .A1(n526), .A2(n657), .ZN(n528) );
  INV_X1 U616 ( .A(KEYINPUT40), .ZN(n527) );
  XNOR2_X2 U617 ( .A(n528), .B(n527), .ZN(n572) );
  XNOR2_X1 U618 ( .A(G131), .B(KEYINPUT127), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n572), .B(n529), .ZN(G33) );
  INV_X1 U620 ( .A(KEYINPUT44), .ZN(n540) );
  AND2_X1 U621 ( .A1(n540), .A2(KEYINPUT66), .ZN(n546) );
  INV_X1 U622 ( .A(n555), .ZN(n678) );
  NAND2_X1 U623 ( .A1(n533), .A2(n532), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n535), .B(n534), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n538), .A2(n350), .ZN(n539) );
  NOR2_X1 U626 ( .A1(n746), .A2(n540), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n545), .B(n544), .ZN(n553) );
  INV_X1 U629 ( .A(KEYINPUT66), .ZN(n547) );
  OR2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U631 ( .A1(n551), .A2(KEYINPUT66), .ZN(n552) );
  NAND2_X1 U632 ( .A1(n553), .A2(n552), .ZN(n567) );
  NOR2_X1 U633 ( .A1(n555), .A2(n682), .ZN(n556) );
  NAND2_X1 U634 ( .A1(n530), .A2(n556), .ZN(n687) );
  OR2_X1 U635 ( .A1(n554), .A2(n687), .ZN(n558) );
  INV_X1 U636 ( .A(KEYINPUT31), .ZN(n557) );
  XNOR2_X1 U637 ( .A(n558), .B(n557), .ZN(n661) );
  NAND2_X1 U638 ( .A1(n559), .A2(n682), .ZN(n560) );
  OR2_X1 U639 ( .A1(n554), .A2(n560), .ZN(n649) );
  NAND2_X1 U640 ( .A1(n661), .A2(n649), .ZN(n563) );
  INV_X1 U641 ( .A(n672), .ZN(n562) );
  NAND2_X1 U642 ( .A1(n563), .A2(n562), .ZN(n564) );
  AND2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U644 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n570) );
  INV_X1 U645 ( .A(n572), .ZN(n583) );
  INV_X1 U646 ( .A(n573), .ZN(n668) );
  NAND2_X1 U647 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U648 ( .A1(n671), .A2(n670), .ZN(n574) );
  XNOR2_X1 U649 ( .A(n574), .B(KEYINPUT41), .ZN(n698) );
  OR2_X1 U650 ( .A1(n682), .A2(n575), .ZN(n577) );
  INV_X1 U651 ( .A(KEYINPUT28), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n577), .B(n576), .ZN(n580) );
  INV_X1 U653 ( .A(n578), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n596) );
  NOR2_X1 U655 ( .A1(n698), .A2(n596), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT42), .ZN(n747) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n585) );
  INV_X1 U658 ( .A(KEYINPUT46), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n585), .B(n584), .ZN(n612) );
  XNOR2_X1 U660 ( .A(n586), .B(KEYINPUT109), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U662 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n589) );
  XNOR2_X1 U663 ( .A(n590), .B(n589), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n591), .A2(n530), .ZN(n593) );
  INV_X1 U665 ( .A(KEYINPUT110), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n593), .B(n592), .ZN(n743) );
  INV_X1 U667 ( .A(n743), .ZN(n601) );
  XNOR2_X1 U668 ( .A(KEYINPUT47), .B(KEYINPUT70), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT76), .ZN(n599) );
  INV_X1 U670 ( .A(n596), .ZN(n598) );
  AND2_X1 U671 ( .A1(n598), .A2(n597), .ZN(n656) );
  NAND2_X1 U672 ( .A1(n599), .A2(n656), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n352), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n672), .A2(KEYINPUT47), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT81), .ZN(n607) );
  INV_X1 U677 ( .A(n656), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n605), .A2(KEYINPUT47), .ZN(n606) );
  AND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT83), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n614) );
  INV_X1 U683 ( .A(KEYINPUT48), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n614), .B(n613), .ZN(n618) );
  AND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  AND2_X2 U686 ( .A1(n618), .A2(n617), .ZN(n734) );
  NAND2_X1 U687 ( .A1(n665), .A2(KEYINPUT2), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n704) );
  INV_X2 U689 ( .A(n704), .ZN(n714) );
  NAND2_X1 U690 ( .A1(n714), .A2(G475), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT59), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(n626) );
  INV_X1 U693 ( .A(G952), .ZN(n625) );
  NOR2_X2 U694 ( .A1(n626), .A2(n718), .ZN(n627) );
  XNOR2_X1 U695 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U696 ( .A1(n714), .A2(G217), .ZN(n630) );
  XNOR2_X1 U697 ( .A(n628), .B(KEYINPUT121), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X2 U699 ( .A1(n631), .A2(n718), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n632), .B(KEYINPUT122), .ZN(G66) );
  NAND2_X1 U701 ( .A1(n714), .A2(G210), .ZN(n637) );
  XNOR2_X1 U702 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n634), .B(KEYINPUT55), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n633), .B(n635), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X2 U706 ( .A1(n638), .A2(n718), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U708 ( .A1(n704), .A2(n640), .ZN(n644) );
  XNOR2_X1 U709 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U711 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n645), .A2(n718), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n647), .B(n646), .ZN(G57) );
  NOR2_X1 U715 ( .A1(n649), .A2(n659), .ZN(n648) );
  XOR2_X1 U716 ( .A(G104), .B(n648), .Z(G6) );
  NOR2_X1 U717 ( .A1(n649), .A2(n662), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U720 ( .A(G107), .B(n652), .ZN(G9) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n655) );
  INV_X1 U722 ( .A(n662), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n653), .A2(n656), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G30) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(G146), .ZN(G48) );
  NOR2_X1 U727 ( .A1(n659), .A2(n661), .ZN(n660) );
  XOR2_X1 U728 ( .A(G113), .B(n660), .Z(G15) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n664) );
  XNOR2_X1 U730 ( .A(G116), .B(KEYINPUT113), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(G18) );
  XOR2_X1 U732 ( .A(n665), .B(KEYINPUT2), .Z(n666) );
  NOR2_X1 U733 ( .A1(n666), .A2(G953), .ZN(n702) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U739 ( .A(KEYINPUT117), .B(n677), .Z(n693) );
  NOR2_X1 U740 ( .A1(n678), .A2(n530), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n679), .B(KEYINPUT50), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n680), .A2(n496), .ZN(n681) );
  XOR2_X1 U743 ( .A(KEYINPUT49), .B(n681), .Z(n683) );
  NAND2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U746 ( .A(n686), .B(KEYINPUT115), .ZN(n688) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U748 ( .A(KEYINPUT51), .B(n689), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n698), .A2(n690), .ZN(n691) );
  XNOR2_X1 U750 ( .A(KEYINPUT116), .B(n691), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT118), .ZN(n695) );
  XNOR2_X1 U753 ( .A(KEYINPUT52), .B(n695), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n675), .A2(n698), .ZN(n699) );
  NOR2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT53), .B(n703), .Z(G75) );
  BUF_X1 U759 ( .A(n704), .Z(n706) );
  NOR2_X1 U760 ( .A1(n706), .A2(n705), .ZN(n712) );
  XOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n708) );
  XNOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n710) );
  XOR2_X1 U764 ( .A(n710), .B(n709), .Z(n711) );
  XNOR2_X1 U765 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U766 ( .A1(n718), .A2(n713), .ZN(G54) );
  NAND2_X1 U767 ( .A1(n714), .A2(G478), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n718), .A2(n717), .ZN(G63) );
  NAND2_X1 U770 ( .A1(n719), .A2(n735), .ZN(n724) );
  XOR2_X1 U771 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n721) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U773 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U776 ( .A(KEYINPUT124), .B(n725), .ZN(n730) );
  XOR2_X1 U777 ( .A(n726), .B(G101), .Z(n728) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(G69) );
  XNOR2_X1 U780 ( .A(KEYINPUT125), .B(n731), .ZN(n733) );
  XNOR2_X1 U781 ( .A(n733), .B(n732), .ZN(n738) );
  XOR2_X1 U782 ( .A(n738), .B(n734), .Z(n736) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U784 ( .A(n737), .B(KEYINPUT126), .ZN(n742) );
  XNOR2_X1 U785 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U788 ( .A1(n742), .A2(n741), .ZN(G72) );
  XNOR2_X1 U789 ( .A(KEYINPUT37), .B(KEYINPUT114), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U791 ( .A(G125), .B(n745), .ZN(G27) );
  XOR2_X1 U792 ( .A(G122), .B(n746), .Z(G24) );
  XOR2_X1 U793 ( .A(G137), .B(n747), .Z(G39) );
endmodule

