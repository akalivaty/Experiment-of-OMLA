//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  NOR2_X1   g0019(.A1(new_n209), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT0), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n221), .A2(new_n222), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n219), .B(new_n229), .C1(new_n222), .C2(new_n221), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0031(.A(G226), .B(G232), .Z(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G97), .B(G107), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT71), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n224), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n224), .A2(new_n262), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n259), .B1(new_n260), .B2(new_n261), .C1(new_n202), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n223), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT11), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n264), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n268));
  OR3_X1    g0068(.A1(new_n258), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n253), .A2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n266), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(KEYINPUT77), .A3(new_n254), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT77), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n255), .B2(new_n266), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n276), .A2(G68), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(G232), .A4(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n280), .A2(new_n282), .A3(G226), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G97), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n291), .A2(KEYINPUT72), .A3(new_n292), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G238), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n253), .B(G274), .C1(G41), .C2(G45), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n289), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(KEYINPUT80), .A3(KEYINPUT13), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT80), .A2(KEYINPUT13), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n289), .A2(new_n297), .A3(new_n298), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(G179), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n289), .A2(new_n297), .A3(new_n306), .A4(new_n298), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n304), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT14), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g0110(.A(KEYINPUT14), .B(new_n304), .C1(new_n305), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n279), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n300), .A2(new_n302), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G190), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n307), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n316), .A3(new_n278), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n295), .A2(G244), .A3(new_n296), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n298), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n280), .A2(new_n282), .A3(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT3), .B(G33), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT73), .A3(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(G238), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n280), .A2(new_n282), .A3(G232), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n280), .A2(new_n282), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(new_n284), .B1(G107), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n288), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n319), .A2(new_n333), .A3(new_n298), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n321), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n336));
  AOI22_X1  g0136(.A1(KEYINPUT75), .A2(new_n320), .B1(new_n331), .B2(new_n288), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT76), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n334), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  OR2_X1    g0141(.A1(KEYINPUT78), .A2(G200), .ZN(new_n342));
  NAND2_X1  g0142(.A1(KEYINPUT78), .A2(G200), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n336), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT8), .B(G58), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(G20), .B2(G77), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT15), .B(G87), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n350), .B1(new_n260), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n266), .B1(new_n261), .B2(new_n255), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n276), .A2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n341), .A2(new_n346), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n340), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n336), .A2(new_n339), .A3(new_n304), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n318), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n255), .A2(new_n266), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(G50), .A3(new_n270), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n347), .A2(new_n260), .B1(new_n365), .B2(new_n263), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G20), .B2(new_n203), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n364), .B1(G50), .B2(new_n254), .C1(new_n367), .C2(new_n272), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(KEYINPUT9), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(KEYINPUT9), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n329), .A2(G1698), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(G222), .B1(G77), .B2(new_n329), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n324), .A2(new_n326), .A3(G223), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n291), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n295), .A2(G226), .A3(new_n296), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n298), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n369), .A2(new_n370), .B1(G190), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n345), .B1(new_n374), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT79), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT10), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(KEYINPUT10), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n378), .A2(new_n381), .A3(KEYINPUT10), .A4(new_n379), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT84), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n291), .A2(G232), .A3(new_n292), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n298), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n280), .A2(new_n282), .A3(G226), .A4(G1698), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n280), .A2(new_n282), .A3(G223), .A4(new_n284), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI211_X1 g0193(.A(G190), .B(new_n389), .C1(new_n288), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n288), .ZN(new_n395));
  INV_X1    g0195(.A(new_n389), .ZN(new_n396));
  AOI21_X1  g0196(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n387), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n393), .B2(new_n288), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(KEYINPUT84), .C1(G200), .C2(new_n399), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n347), .A2(new_n271), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n404), .A2(new_n272), .B1(new_n255), .B2(new_n347), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT16), .ZN(new_n407));
  INV_X1    g0207(.A(G159), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT81), .B1(new_n263), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT81), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n349), .A2(new_n410), .A3(G159), .ZN(new_n411));
  XNOR2_X1  g0211(.A(G58), .B(G68), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n409), .A2(new_n411), .B1(new_n412), .B2(G20), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT82), .B1(new_n281), .B2(G33), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT82), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(new_n262), .A3(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n416), .A3(new_n282), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n325), .B2(G20), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n256), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n413), .B1(new_n422), .B2(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n329), .A2(new_n224), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n424), .A2(new_n418), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT83), .ZN(new_n426));
  NOR3_X1   g0226(.A1(new_n425), .A2(new_n426), .A3(new_n256), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n407), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n329), .B2(new_n224), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n418), .B(G20), .C1(new_n280), .C2(new_n282), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT16), .A3(new_n413), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n432), .A2(new_n266), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n406), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n403), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n403), .B2(new_n434), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n399), .A2(G179), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n399), .A2(new_n304), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n439), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n432), .A2(new_n266), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n426), .B1(new_n425), .B2(new_n256), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n413), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n448), .B2(new_n407), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT18), .B(new_n444), .C1(new_n449), .C2(new_n406), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n438), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n368), .B1(new_n377), .B2(G169), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n377), .A2(new_n358), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR4_X1   g0260(.A1(new_n362), .A2(new_n386), .A3(new_n453), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n462), .A2(new_n212), .A3(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n465), .A2(new_n224), .B1(new_n261), .B2(new_n263), .ZN(new_n466));
  INV_X1    g0266(.A(G107), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n420), .B2(new_n421), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n266), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(G33), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT86), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n363), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n255), .A2(new_n212), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT85), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G41), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n253), .B(G45), .C1(new_n478), .C2(KEYINPUT5), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n288), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n253), .A2(G45), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(G274), .A4(new_n481), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(G1698), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(new_n284), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n325), .A2(new_n495), .A3(G244), .A4(new_n284), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n288), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(new_n496), .ZN(new_n500));
  INV_X1    g0300(.A(new_n492), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n500), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n489), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n477), .B1(new_n503), .B2(G200), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT88), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n503), .B2(new_n400), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n291), .B1(new_n507), .B2(KEYINPUT87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n497), .A2(new_n498), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n488), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(KEYINPUT88), .A3(G190), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n358), .B(new_n489), .C1(new_n499), .C2(new_n502), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n477), .C1(new_n510), .C2(G169), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(new_n284), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G294), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n322), .C2(new_n213), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n288), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n482), .A2(G264), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n487), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  XOR2_X1   g0321(.A(KEYINPUT92), .B(KEYINPUT22), .Z(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(new_n224), .A3(G87), .A4(new_n325), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n260), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(G20), .B2(new_n467), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n224), .A2(KEYINPUT23), .A3(G107), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n280), .A2(new_n282), .A3(new_n224), .A4(G87), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT92), .B(KEYINPUT22), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n523), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n523), .A2(new_n529), .A3(KEYINPUT24), .A4(new_n532), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n266), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT25), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n254), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n255), .A2(KEYINPUT25), .A3(new_n467), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n473), .A2(G107), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n517), .A2(new_n288), .B1(new_n482), .B2(G264), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(G190), .A3(new_n487), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n521), .A2(new_n537), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  OR2_X1    g0344(.A1(new_n472), .A2(new_n351), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n224), .B1(new_n286), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G87), .B2(new_n206), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n280), .A2(new_n282), .A3(new_n224), .A4(G68), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n260), .B2(new_n212), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(new_n266), .B1(new_n255), .B2(new_n351), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G116), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n280), .A2(new_n282), .A3(G238), .A4(new_n284), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(KEYINPUT89), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(KEYINPUT89), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n288), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n484), .A2(G250), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(new_n291), .B1(new_n485), .B2(G274), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n358), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n561), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(KEYINPUT89), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n325), .A2(new_n565), .A3(G238), .A4(new_n284), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n564), .A2(new_n566), .A3(new_n554), .A4(new_n555), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n567), .B2(new_n288), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n553), .B(new_n562), .C1(G169), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n551), .A2(new_n266), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n351), .A2(new_n255), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n471), .A2(new_n363), .A3(G87), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n559), .A2(G190), .A3(new_n561), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n344), .C2(new_n568), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n544), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n512), .A2(new_n514), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT91), .ZN(new_n578));
  INV_X1    g0378(.A(new_n481), .ZN(new_n579));
  OAI211_X1 g0379(.A(G270), .B(new_n291), .C1(new_n579), .C2(new_n479), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n487), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(new_n284), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT90), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT90), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n325), .A2(new_n584), .A3(G257), .A4(new_n284), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n325), .A2(G264), .A3(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n329), .A2(G303), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n581), .B1(new_n588), .B2(new_n288), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G179), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n592));
  OAI21_X1  g0392(.A(G116), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n275), .B2(new_n273), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n265), .A2(new_n223), .B1(G20), .B2(new_n524), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n491), .B(new_n224), .C1(G33), .C2(new_n212), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT20), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(G116), .B2(new_n254), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n578), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  AOI211_X1 g0401(.A(new_n358), .B(new_n581), .C1(new_n588), .C2(new_n288), .ZN(new_n602));
  INV_X1    g0402(.A(new_n598), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(KEYINPUT20), .A3(new_n596), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n604), .B1(new_n524), .B2(new_n255), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n273), .A2(new_n275), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G116), .A3(new_n471), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(KEYINPUT91), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n537), .A2(new_n541), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n520), .A2(G169), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT93), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(new_n358), .B2(new_n520), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n304), .B1(new_n542), .B2(new_n487), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(KEYINPUT93), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n611), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  OAI21_X1  g0418(.A(G169), .B1(new_n594), .B2(new_n599), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n589), .ZN(new_n620));
  INV_X1    g0420(.A(new_n589), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n608), .A3(KEYINPUT21), .A4(G169), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n621), .A2(new_n400), .ZN(new_n624));
  INV_X1    g0424(.A(G200), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n600), .B1(new_n625), .B2(new_n589), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n610), .A2(new_n617), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n577), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n461), .A2(new_n629), .ZN(G372));
  NAND3_X1  g0430(.A1(new_n610), .A2(new_n617), .A3(new_n623), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n514), .A3(new_n512), .A4(new_n576), .ZN(new_n632));
  INV_X1    g0432(.A(new_n569), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n559), .A2(new_n561), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n304), .B1(new_n545), .B2(new_n552), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n634), .B2(new_n345), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n562), .A2(new_n635), .B1(new_n637), .B2(new_n574), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n474), .A2(new_n476), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n503), .A2(new_n304), .B1(new_n639), .B2(new_n469), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(KEYINPUT26), .A3(new_n513), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n569), .A2(new_n575), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n514), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n633), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT94), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n632), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AOI211_X1 g0447(.A(KEYINPUT94), .B(new_n633), .C1(new_n641), .C2(new_n644), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n461), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n428), .A2(new_n433), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n405), .A3(new_n398), .A4(new_n402), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n403), .A2(new_n434), .A3(new_n435), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n317), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n312), .B2(new_n361), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT95), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n409), .A2(new_n411), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n412), .A2(G20), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n420), .A2(new_n421), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G68), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n426), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT16), .B1(new_n664), .B2(new_n447), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n405), .B1(new_n665), .B2(new_n445), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT18), .B1(new_n666), .B2(new_n444), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n434), .A2(new_n439), .A3(new_n442), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n658), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n443), .A2(KEYINPUT95), .A3(new_n450), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n384), .B(new_n385), .C1(new_n657), .C2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(new_n459), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n650), .A2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(G13), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n253), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI211_X1 g0483(.A(new_n600), .B(new_n683), .C1(new_n610), .C2(new_n623), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n601), .A2(new_n620), .A3(new_n609), .A4(new_n622), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n608), .B2(new_n682), .ZN(new_n686));
  OAI211_X1 g0486(.A(G330), .B(new_n627), .C1(new_n684), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n611), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n617), .B(new_n544), .C1(new_n689), .C2(new_n683), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n520), .A2(new_n358), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n615), .B2(KEYINPUT93), .ZN(new_n692));
  INV_X1    g0492(.A(new_n616), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n682), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n685), .A2(new_n683), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n685), .A2(new_n617), .A3(new_n544), .A4(new_n683), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n694), .A2(new_n683), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT96), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n220), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n227), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n649), .A2(new_n683), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n632), .A2(new_n645), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n683), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n713), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n512), .A2(new_n514), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n624), .A2(new_n626), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n694), .A2(new_n685), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(new_n722), .A3(new_n576), .A4(new_n683), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n503), .A2(new_n590), .ZN(new_n724));
  AND4_X1   g0524(.A1(KEYINPUT97), .A2(new_n542), .A3(new_n559), .A4(new_n561), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT97), .B1(new_n568), .B2(new_n542), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n727), .A3(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n542), .A2(new_n559), .A3(new_n561), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT97), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n568), .A2(KEYINPUT97), .A3(new_n542), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n507), .A2(KEYINPUT87), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n288), .A3(new_n509), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(new_n489), .A3(new_n602), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n729), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT98), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n589), .A2(G179), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n503), .A2(new_n634), .A3(new_n520), .A4(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n728), .A2(new_n738), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n728), .A2(new_n738), .A3(new_n741), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n683), .B1(new_n743), .B2(KEYINPUT98), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n723), .A2(KEYINPUT31), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n719), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n711), .B1(new_n749), .B2(G1), .ZN(G364));
  NAND2_X1  g0550(.A1(new_n676), .A2(G45), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT99), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n253), .B1(new_n751), .B2(KEYINPUT99), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n706), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n627), .B1(new_n684), .B2(new_n686), .ZN(new_n757));
  INV_X1    g0557(.A(G330), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n756), .B1(new_n759), .B2(new_n688), .ZN(new_n760));
  OR3_X1    g0560(.A1(KEYINPUT100), .A2(G13), .A3(G33), .ZN(new_n761));
  OAI21_X1  g0561(.A(KEYINPUT100), .B1(G13), .B2(G33), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n223), .B1(G20), .B2(new_n304), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n705), .A2(new_n325), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n227), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G45), .B2(new_n251), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n705), .A2(new_n329), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G355), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G116), .B2(new_n220), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n767), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n400), .A2(G20), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n344), .A2(G179), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n224), .A2(new_n400), .A3(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n345), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n224), .A2(new_n400), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n358), .A2(new_n625), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G326), .ZN(new_n787));
  INV_X1    g0587(.A(new_n775), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n784), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI22_X1  g0590(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n775), .A2(new_n358), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G329), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n793), .A2(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n224), .B1(new_n795), .B2(G190), .ZN(new_n799));
  INV_X1    g0599(.A(G294), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n783), .A2(G179), .A3(new_n625), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n329), .B1(new_n799), .B2(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n782), .A2(new_n791), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n780), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G87), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n806), .B(new_n325), .C1(new_n467), .C2(new_n777), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  INV_X1    g0608(.A(new_n801), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n809), .A2(G58), .B1(new_n785), .B2(G50), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n810), .B1(new_n256), .B2(new_n789), .C1(new_n261), .C2(new_n793), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n796), .A2(KEYINPUT32), .A3(new_n408), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n796), .B2(new_n408), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n212), .B2(new_n799), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n804), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n766), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n774), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n757), .B2(new_n765), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n760), .B1(new_n756), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT102), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND3_X1  g0622(.A1(new_n359), .A2(new_n360), .A3(new_n683), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n355), .B1(new_n340), .B2(G190), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(new_n346), .B1(new_n355), .B2(new_n682), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n359), .A2(new_n360), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n712), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n338), .B1(new_n337), .B2(new_n334), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n358), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g0631(.A1(new_n355), .A2(new_n831), .A3(new_n360), .A4(new_n683), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n355), .A2(new_n682), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n357), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n834), .B2(new_n361), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n683), .B(new_n835), .C1(new_n647), .C2(new_n648), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n755), .B1(new_n837), .B2(new_n748), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n748), .B2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n763), .A2(new_n766), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n756), .B1(new_n261), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n776), .A2(G87), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n467), .B2(new_n780), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n786), .A2(new_n781), .B1(new_n801), .B2(new_n800), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n793), .A2(new_n524), .B1(new_n796), .B2(new_n794), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n329), .B1(new_n799), .B2(new_n212), .C1(new_n789), .C2(new_n778), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G58), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n325), .B1(new_n799), .B2(new_n848), .C1(new_n796), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n776), .A2(G68), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n202), .B2(new_n780), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n365), .A2(new_n789), .B1(new_n801), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n793), .A2(new_n408), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(G137), .C2(new_n785), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n850), .B(new_n852), .C1(new_n856), .C2(KEYINPUT34), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n847), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n841), .B1(new_n817), .B2(new_n859), .C1(new_n835), .C2(new_n764), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n839), .A2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n676), .A2(new_n253), .ZN(new_n862));
  NOR2_X1   g0662(.A1(KEYINPUT105), .A2(KEYINPUT16), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n431), .A2(new_n413), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n256), .B1(new_n421), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n863), .B1(new_n867), .B2(new_n661), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n868), .A3(new_n266), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n405), .ZN(new_n870));
  INV_X1    g0670(.A(new_n680), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n438), .B2(new_n451), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n442), .A2(new_n680), .B1(new_n869), .B2(new_n405), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n434), .B2(new_n403), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n870), .B1(new_n444), .B2(new_n871), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n652), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(KEYINPUT106), .A3(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n444), .B1(new_n449), .B2(new_n406), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n871), .B1(new_n449), .B2(new_n406), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(new_n652), .A4(new_n878), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n879), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n874), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n874), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n874), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n669), .A2(new_n655), .A3(new_n670), .ZN(new_n892));
  INV_X1    g0692(.A(new_n884), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n883), .A2(new_n884), .A3(new_n652), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT37), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n892), .A2(new_n893), .B1(new_n885), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n890), .B(new_n891), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n312), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n683), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n900), .A2(new_n903), .B1(new_n671), .B2(new_n680), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n279), .A2(new_n682), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n312), .A2(new_n317), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n279), .B(new_n682), .C1(new_n310), .C2(new_n311), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT103), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n836), .B2(new_n823), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n874), .A2(new_n886), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n891), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n913), .B2(new_n914), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n904), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n714), .A2(new_n461), .A3(new_n718), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n673), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n921), .B(new_n923), .Z(new_n924));
  NAND2_X1  g0724(.A1(new_n895), .A2(new_n885), .ZN(new_n925));
  INV_X1    g0725(.A(new_n670), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT95), .B1(new_n443), .B2(new_n450), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n926), .A2(new_n438), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n925), .B1(new_n928), .B2(new_n884), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n443), .A2(new_n450), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n872), .B1(new_n655), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT106), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n932));
  AND4_X1   g0732(.A1(new_n878), .A2(new_n883), .A3(new_n884), .A4(new_n652), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(new_n882), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n929), .A2(new_n897), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n742), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT31), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n629), .B2(new_n683), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n743), .A2(KEYINPUT98), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n940), .A2(new_n682), .A3(new_n742), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n937), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n827), .B1(new_n909), .B2(new_n911), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT40), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n919), .A2(new_n946), .A3(new_n942), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(G330), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n461), .A2(G330), .A3(new_n942), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n461), .A2(new_n942), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n862), .B1(new_n924), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n952), .B2(new_n924), .ZN(new_n954));
  INV_X1    g0754(.A(new_n465), .ZN(new_n955));
  OAI211_X1 g0755(.A(G116), .B(new_n225), .C1(new_n955), .C2(KEYINPUT35), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(KEYINPUT35), .B2(new_n955), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT36), .Z(new_n958));
  OAI21_X1  g0758(.A(G77), .B1(new_n848), .B2(new_n256), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n227), .A2(new_n959), .B1(G50), .B2(new_n256), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n675), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(G367));
  NAND2_X1  g0762(.A1(new_n477), .A2(new_n682), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n512), .A2(new_n514), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n640), .A2(new_n513), .A3(new_n682), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(new_n699), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT42), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n720), .A2(new_n694), .A3(new_n963), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n682), .B1(new_n969), .B2(new_n514), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n967), .B2(KEYINPUT42), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n573), .A2(new_n683), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n633), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n643), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n968), .A2(new_n971), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT108), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT108), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n968), .A2(new_n971), .A3(new_n978), .A4(new_n975), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n968), .A2(new_n971), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n974), .B(KEYINPUT43), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n981), .B1(new_n980), .B2(new_n984), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(new_n698), .B2(new_n966), .ZN(new_n988));
  INV_X1    g0788(.A(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n698), .A2(new_n966), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(new_n985), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n706), .B(KEYINPUT41), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n701), .B(KEYINPUT96), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n966), .ZN(new_n996));
  INV_X1    g0796(.A(new_n966), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n703), .B2(new_n997), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n995), .A2(KEYINPUT44), .A3(new_n966), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n999), .A2(new_n1003), .A3(new_n698), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n698), .B1(new_n999), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n697), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n699), .B1(new_n687), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n687), .B2(new_n1007), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT29), .B1(new_n649), .B2(new_n683), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n748), .B(new_n1009), .C1(new_n1010), .C2(new_n717), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT110), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n719), .A2(new_n1013), .A3(new_n748), .A4(new_n1009), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1006), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n993), .B1(new_n1015), .B2(new_n749), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n988), .B(new_n991), .C1(new_n1016), .C2(new_n754), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n240), .A2(new_n705), .A3(new_n325), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n767), .B1(new_n220), .B2(new_n351), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n755), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n799), .A2(new_n256), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n805), .B2(G58), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n796), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n329), .B1(new_n1023), .B2(G137), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(new_n261), .C2(new_n777), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n809), .A2(G150), .B1(G50), .B2(new_n792), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n853), .B2(new_n786), .C1(new_n408), .C2(new_n789), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n780), .B2(new_n524), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1023), .A2(G317), .B1(new_n785), .B2(G311), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n789), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(G294), .B1(G283), .B2(new_n792), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n325), .B1(new_n809), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n467), .B2(new_n799), .C1(new_n777), .C2(new_n212), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1025), .A2(new_n1027), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT47), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n817), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1020), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n765), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n974), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1017), .A2(new_n1043), .ZN(G387));
  AOI22_X1  g0844(.A1(new_n785), .A2(G322), .B1(new_n792), .B2(G303), .ZN(new_n1045));
  INV_X1    g0845(.A(G317), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(new_n794), .B2(new_n789), .C1(new_n1046), .C2(new_n801), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n778), .B2(new_n799), .C1(new_n800), .C2(new_n780), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n329), .B1(new_n787), .B2(new_n796), .C1(new_n777), .C2(new_n524), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n805), .A2(G77), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n365), .B2(new_n796), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT112), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n348), .A2(new_n1032), .B1(new_n809), .B2(G50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n408), .B2(new_n786), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n799), .A2(new_n351), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n325), .B1(new_n256), .B2(new_n793), .C1(new_n777), .C2(new_n212), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT113), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n817), .B1(new_n1054), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n708), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n771), .A2(new_n1065), .B1(new_n467), .B2(new_n705), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT111), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT111), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n236), .A2(G45), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT50), .B1(new_n347), .B2(G50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n708), .A3(new_n1071), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n347), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n768), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1067), .B(new_n1068), .C1(new_n1069), .C2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n756), .B(new_n1064), .C1(new_n767), .C2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n690), .A2(new_n695), .A3(new_n765), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1076), .A2(new_n1077), .B1(new_n754), .B2(new_n1009), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n749), .A2(new_n1009), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1011), .A2(new_n706), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1006), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1011), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n706), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n706), .A4(new_n1084), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1006), .A2(new_n754), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n793), .A2(new_n800), .B1(new_n796), .B2(new_n802), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n325), .B(new_n1089), .C1(G303), .C2(new_n1032), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n777), .A2(new_n467), .B1(new_n778), .B2(new_n780), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n799), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(G116), .B2(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n786), .A2(new_n1046), .B1(new_n801), .B2(new_n794), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT52), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1090), .A2(new_n1093), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n789), .A2(new_n202), .B1(new_n796), .B2(new_n853), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n329), .B(new_n1099), .C1(new_n348), .C2(new_n792), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n842), .B1(new_n256), .B2(new_n780), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n799), .A2(new_n261), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n786), .A2(new_n365), .B1(new_n801), .B2(new_n408), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT51), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1100), .A2(new_n1103), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n817), .B1(new_n1098), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n246), .A2(new_n768), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n766), .B(new_n765), .C1(new_n705), .C2(G97), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n756), .B(new_n1109), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n997), .B2(new_n1042), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1113), .ZN(G390));
  NAND3_X1  g0914(.A1(new_n942), .A2(new_n943), .A3(G330), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT115), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n942), .A2(new_n943), .A3(new_n1117), .A4(G330), .ZN(new_n1118));
  OAI211_X1 g0918(.A(G330), .B(new_n835), .C1(new_n745), .C2(new_n746), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n912), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n836), .A2(new_n823), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1119), .A2(new_n912), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n825), .A2(new_n826), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n823), .B1(new_n716), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n942), .A2(G330), .A3(new_n835), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n912), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n922), .A2(new_n673), .A3(new_n950), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n909), .A2(new_n911), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n891), .B1(new_n896), .B2(new_n898), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n902), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n903), .B1(new_n1122), .B2(new_n1134), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n900), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1124), .B(new_n1137), .C1(new_n1138), .C2(new_n900), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n706), .B1(new_n1133), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT116), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1142), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT118), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1130), .A2(new_n1149), .A3(new_n1132), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1121), .A2(new_n1122), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1151));
  OAI21_X1  g0951(.A(KEYINPUT118), .B1(new_n1151), .B2(new_n1131), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT116), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n706), .C1(new_n1133), .C2(new_n1143), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1145), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n754), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1143), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n889), .A2(new_n899), .A3(new_n763), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n840), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n755), .B1(new_n348), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n325), .B1(new_n1163), .B2(new_n796), .C1(new_n777), .C2(new_n202), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G159), .B2(new_n1092), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n780), .A2(new_n365), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT53), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G137), .A2(new_n1032), .B1(new_n809), .B2(G132), .ZN(new_n1168));
  XOR2_X1   g0968(.A(KEYINPUT54), .B(G143), .Z(new_n1169));
  AOI22_X1  g0969(.A1(new_n785), .A2(G128), .B1(new_n792), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n806), .A2(new_n329), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT119), .Z(new_n1173));
  OAI22_X1  g0973(.A1(new_n800), .A2(new_n796), .B1(new_n801), .B2(new_n524), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G97), .B2(new_n792), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1102), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1032), .A2(G107), .B1(new_n785), .B2(G283), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n851), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1171), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1162), .B1(new_n1179), .B2(new_n766), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1159), .B1(new_n1160), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1157), .A2(new_n1181), .ZN(G378));
  NAND2_X1  g0982(.A1(new_n368), .A2(new_n871), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n386), .B2(new_n460), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n384), .A2(new_n459), .A3(new_n385), .A4(new_n1183), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n948), .B2(G330), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n758), .B(new_n1190), .C1(new_n945), .C2(new_n947), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n921), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1136), .A2(new_n942), .A3(new_n943), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n942), .A2(new_n943), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT40), .B1(new_n918), .B2(new_n891), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1195), .A2(KEYINPUT40), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1190), .B1(new_n1198), .B2(new_n758), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n915), .A2(new_n920), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n946), .B1(new_n1196), .B2(new_n1136), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n946), .B1(new_n887), .B2(new_n888), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(new_n944), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G330), .B(new_n1191), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n904), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1132), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1206), .A2(KEYINPUT57), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1209));
  OR3_X1    g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n707), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n754), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT123), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1190), .A2(new_n763), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G33), .A2(G41), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT120), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G50), .B(new_n1215), .C1(new_n478), .C2(new_n329), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n786), .A2(new_n524), .B1(new_n789), .B2(new_n212), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n793), .A2(new_n351), .B1(new_n796), .B2(new_n778), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n478), .B(new_n329), .C1(new_n801), .C2(new_n467), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n1021), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n776), .A2(G58), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1055), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT58), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1216), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1032), .A2(G132), .B1(G137), .B2(new_n792), .ZN(new_n1226));
  INV_X1    g1026(.A(G128), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(new_n801), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n785), .A2(G125), .B1(new_n1092), .B2(G150), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT121), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n805), .C2(new_n1169), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT59), .Z(new_n1232));
  OR2_X1    g1032(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1023), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n1215), .C1(new_n777), .C2(new_n408), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1225), .B1(new_n1224), .B2(new_n1223), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n766), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n756), .B1(new_n202), .B2(new_n840), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1213), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1211), .A2(new_n1212), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1158), .B1(new_n1194), .B2(new_n1205), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1240), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT123), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1210), .A2(new_n1245), .ZN(G375));
  NAND3_X1  g1046(.A1(new_n1123), .A2(new_n1131), .A3(new_n1129), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1153), .A2(new_n992), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1222), .B(new_n325), .C1(new_n1227), .C2(new_n796), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n780), .A2(new_n408), .B1(new_n202), .B2(new_n799), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n809), .A2(G137), .B1(new_n785), .B2(G132), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1032), .A2(new_n1169), .B1(new_n792), .B2(G150), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n329), .B1(new_n467), .B2(new_n793), .C1(new_n777), .C2(new_n261), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n780), .A2(new_n212), .B1(new_n351), .B2(new_n799), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n789), .A2(new_n524), .B1(new_n796), .B2(new_n781), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n786), .A2(new_n800), .B1(new_n801), .B2(new_n778), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n766), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n755), .C1(G68), .C2(new_n1161), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT124), .Z(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n912), .B2(new_n763), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n1130), .B2(new_n754), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1248), .A2(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(new_n1181), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(KEYINPUT116), .A2(new_n1144), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1156), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1210), .A2(new_n1245), .A3(new_n1268), .ZN(new_n1269));
  OR4_X1    g1069(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1270));
  OR4_X1    g1070(.A1(G387), .A2(new_n1269), .A3(G381), .A4(new_n1270), .ZN(G407));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(G343), .C2(new_n1269), .ZN(G409));
  NOR3_X1   g1072(.A1(new_n1208), .A2(new_n1209), .A3(new_n707), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1274));
  OAI21_X1  g1074(.A(G378), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1206), .A2(new_n992), .A3(new_n1207), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(new_n1240), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1194), .B2(new_n1205), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1194), .A2(new_n1205), .A3(new_n1281), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n754), .A3(new_n1284), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1157), .A3(new_n1285), .A4(new_n1181), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1247), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1288), .A2(new_n706), .A3(new_n1133), .A4(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(G384), .A3(new_n1264), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1290), .B2(new_n1264), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1275), .A2(new_n1278), .A3(new_n1286), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT126), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1277), .A2(G2897), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1290), .A2(new_n1264), .ZN(new_n1302));
  INV_X1    g1102(.A(G384), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1291), .A3(new_n1299), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1194), .A2(new_n1281), .A3(new_n1205), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1307), .A2(new_n1282), .A3(new_n1158), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1279), .A2(new_n1240), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1277), .B1(new_n1310), .B2(new_n1268), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1306), .B1(new_n1311), .B2(new_n1275), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(G393), .B(new_n821), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(G390), .A2(new_n1043), .A3(new_n1017), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1017), .B2(new_n1043), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1314), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G390), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1312), .A2(KEYINPUT61), .A3(new_n1322), .ZN(new_n1323));
  OR2_X1    g1123(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1295), .A2(new_n1325), .A3(new_n1296), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1298), .A2(new_n1323), .A3(new_n1324), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1311), .A2(new_n1275), .A3(new_n1330), .A4(new_n1294), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1306), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1268), .B1(new_n1210), .B2(new_n1245), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1286), .A2(new_n1278), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1328), .A2(new_n1329), .A3(new_n1331), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1322), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1327), .A2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1269), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1339), .B1(new_n1340), .B2(new_n1333), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1339), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1269), .B(new_n1275), .C1(new_n1342), .C2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1341), .A2(new_n1344), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1322), .ZN(G402));
endmodule


