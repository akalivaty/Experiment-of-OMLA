//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1191,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n463), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n464), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(KEYINPUT67), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n464), .A2(G138), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n465), .C1(new_n461), .C2(new_n462), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n483), .B1(new_n487), .B2(new_n484), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n476), .B2(G126), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT69), .A2(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT69), .A2(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT5), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(KEYINPUT5), .C1(new_n497), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n496), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n506), .B1(new_n500), .B2(new_n502), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(G88), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n513), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n515), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT6), .B(G651), .Z(new_n523));
  AOI211_X1 g098(.A(new_n523), .B(new_n506), .C1(new_n500), .C2(new_n502), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n517), .A2(G51), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n525), .A2(new_n526), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n524), .A2(G90), .B1(G52), .B2(new_n517), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n508), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n512), .A2(G81), .A3(new_n513), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(G43), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n542), .A2(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n512), .A2(G91), .A3(new_n513), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n513), .A2(G543), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n558), .B(new_n562), .C1(new_n563), .C2(new_n534), .ZN(G299));
  NAND2_X1  g139(.A1(new_n524), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n517), .A2(G49), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n534), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G48), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n512), .A2(new_n513), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n570), .A2(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(G72), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G60), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n508), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n534), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT77), .B(new_n576), .C1(new_n508), .C2(new_n577), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n524), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NOR2_X1   g160(.A1(G301), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT69), .B(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n501), .B1(new_n587), .B2(KEYINPUT5), .ZN(new_n588));
  INV_X1    g163(.A(new_n502), .ZN(new_n589));
  OAI211_X1 g164(.A(G66), .B(new_n507), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n503), .A2(G92), .A3(new_n507), .A4(new_n513), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n513), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(KEYINPUT78), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT78), .B1(new_n593), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n586), .B1(new_n602), .B2(new_n585), .ZN(G284));
  AOI21_X1  g178(.A(new_n586), .B1(new_n602), .B2(new_n585), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n512), .A2(G65), .ZN(new_n606));
  NAND2_X1  g181(.A1(G78), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n534), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n558), .A2(new_n562), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n605), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n605), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n602), .B1(new_n613), .B2(G860), .ZN(G148));
  OAI21_X1  g189(.A(new_n613), .B1(new_n599), .B2(new_n600), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n616), .A2(KEYINPUT79), .A3(new_n585), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT79), .B1(new_n616), .B2(new_n585), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n617), .B(new_n618), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g195(.A1(new_n463), .A2(new_n466), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n464), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n476), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n465), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n627), .A2(new_n628), .A3(new_n635), .ZN(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT17), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n652), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n657), .A2(new_n654), .A3(new_n652), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n654), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n653), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n634), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT83), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT85), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n673), .A2(new_n679), .A3(new_n676), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n678), .B(new_n680), .C1(new_n676), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n570), .A2(new_n574), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G16), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT32), .ZN(new_n692));
  OR2_X1    g267(.A1(G6), .A2(G16), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(G1981), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1981), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(G166), .A2(G16), .ZN(new_n703));
  OR2_X1    g278(.A1(G16), .A2(G22), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(G1971), .A3(new_n704), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n689), .B1(new_n702), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n715), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n717), .A2(KEYINPUT34), .A3(new_n701), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n708), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(new_n583), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n580), .B2(new_n581), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n720), .B1(new_n722), .B2(new_n708), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(G1986), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n723), .B(new_n724), .Z(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT87), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n464), .A2(G131), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT88), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n476), .A2(G119), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n465), .A2(G107), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n725), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT91), .Z(new_n742));
  NAND3_X1  g317(.A1(new_n719), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n552), .A2(G16), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n745));
  OR2_X1    g320(.A1(G16), .A2(G19), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n749));
  OAI21_X1  g324(.A(G1341), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n751), .A2(new_n752), .A3(new_n747), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(G168), .A2(G16), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(KEYINPUT95), .C1(G16), .C2(G21), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n757), .B1(new_n758), .B2(new_n756), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n708), .A2(G5), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G301), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n759), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n708), .A2(G4), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n602), .B2(new_n708), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(G1348), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n708), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n610), .B2(new_n708), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1956), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n480), .A2(G29), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n726), .A2(G35), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(G2090), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(KEYINPUT97), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n780), .A2(new_n781), .B1(new_n763), .B2(new_n762), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n464), .A2(G139), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(G127), .B1(new_n461), .B2(new_n462), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n465), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n787), .A2(new_n790), .A3(new_n726), .ZN(new_n791));
  INV_X1    g366(.A(G2072), .ZN(new_n792));
  NOR2_X1   g367(.A1(G29), .A2(G33), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT24), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G34), .ZN(new_n799));
  AOI21_X1  g374(.A(G29), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n473), .B2(G29), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n726), .A2(G32), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n476), .A2(G129), .ZN(new_n805));
  NAND3_X1  g380(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT26), .Z(new_n807));
  AND3_X1   g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n803), .B1(new_n808), .B2(new_n726), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT27), .B(G1996), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n464), .A2(G140), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n476), .A2(G128), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n465), .A2(G116), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n726), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(G2067), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n803), .B(new_n810), .C1(new_n808), .C2(new_n726), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n818), .A2(new_n820), .A3(new_n822), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n812), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n801), .A2(new_n796), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT30), .B(G28), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n829), .A2(new_n726), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n828), .B(new_n832), .C1(new_n726), .C2(new_n633), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n777), .A2(new_n778), .A3(G2090), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n802), .A2(new_n827), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n726), .A2(G27), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT96), .Z(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G164), .B2(new_n726), .ZN(new_n838));
  INV_X1    g413(.A(G2078), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AND4_X1   g415(.A1(new_n773), .A2(new_n782), .A3(new_n835), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n754), .A2(new_n765), .A3(new_n769), .A4(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n743), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n739), .B1(new_n716), .B2(new_n718), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n742), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n844), .A2(KEYINPUT98), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n845), .A2(new_n742), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n842), .B1(new_n845), .B2(new_n742), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n847), .A2(new_n851), .ZN(G311));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n850), .ZN(G150));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n524), .A2(G93), .B1(G55), .B2(new_n517), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n503), .A2(G67), .A3(new_n507), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n534), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n861), .A2(KEYINPUT99), .A3(new_n534), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n854), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n859), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT99), .B1(new_n861), .B2(new_n534), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT100), .A4(new_n855), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n602), .A2(G559), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n863), .A2(new_n551), .A3(new_n866), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n534), .B1(new_n541), .B2(KEYINPUT74), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(KEYINPUT74), .B2(new_n541), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n549), .A2(new_n550), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(new_n865), .A3(new_n855), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n871), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT101), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n879), .B2(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n869), .B1(new_n881), .B2(new_n883), .ZN(G145));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n494), .B(KEYINPUT103), .Z(new_n886));
  NOR2_X1   g461(.A1(new_n787), .A2(new_n790), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n734), .B(new_n623), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n808), .B(new_n817), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n476), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n465), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n464), .A2(new_n895), .A3(G142), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n464), .B2(G142), .ZN(new_n897));
  OAI221_X1 g472(.A(new_n892), .B1(new_n893), .B2(new_n894), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n891), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n890), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n473), .B(KEYINPUT102), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n480), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n633), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n900), .A2(new_n903), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n885), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n905), .A4(new_n904), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(G395));
  XNOR2_X1  g486(.A(new_n690), .B(G288), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n722), .A2(G303), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n722), .A2(G303), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n690), .B(new_n710), .ZN(new_n916));
  NAND2_X1  g491(.A1(G290), .A2(G166), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n722), .A2(G303), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n596), .A2(new_n597), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n517), .A2(G54), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n534), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n610), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(G299), .A2(new_n593), .A3(new_n598), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n610), .B(KEYINPUT105), .C1(new_n923), .C2(new_n926), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n872), .A2(new_n615), .A3(new_n877), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n615), .B1(new_n872), .B2(new_n877), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n878), .A2(new_n616), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n872), .A2(new_n615), .A3(new_n877), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n939), .A2(new_n940), .B1(new_n928), .B2(new_n927), .ZN(new_n941));
  NOR2_X1   g516(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n933), .A2(new_n934), .ZN(new_n945));
  INV_X1    g520(.A(new_n929), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n939), .A3(new_n940), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n927), .A2(new_n928), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n936), .B2(new_n937), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n944), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n922), .B1(new_n943), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n938), .B2(new_n941), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(new_n940), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n950), .B(new_n944), .C1(new_n954), .C2(new_n935), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n921), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n585), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n867), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(G868), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(KEYINPUT107), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n953), .A2(new_n921), .A3(new_n955), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n921), .B1(new_n953), .B2(new_n955), .ZN(new_n963));
  OAI21_X1  g538(.A(G868), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n959), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n960), .A2(new_n966), .ZN(G295));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n965), .ZN(G331));
  AND3_X1   g543(.A1(new_n535), .A2(G286), .A3(new_n536), .ZN(new_n969));
  AOI21_X1  g544(.A(G286), .B1(new_n535), .B2(new_n536), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n872), .A2(new_n877), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n872), .B2(new_n877), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT109), .B1(new_n974), .B2(new_n935), .ZN(new_n975));
  INV_X1    g550(.A(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n878), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n872), .A2(new_n971), .A3(new_n877), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n947), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n949), .A3(new_n978), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n975), .A2(new_n981), .A3(new_n920), .A4(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n928), .A4(new_n932), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n949), .A2(new_n934), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n972), .B2(new_n973), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(new_n982), .A3(KEYINPUT111), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n915), .A2(new_n919), .A3(KEYINPUT110), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n915), .B2(new_n919), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n979), .A2(new_n992), .A3(new_n986), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n983), .A2(new_n994), .A3(new_n905), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n975), .A2(new_n981), .A3(new_n982), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n991), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(new_n905), .A3(new_n983), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n996), .B(KEYINPUT44), .C1(new_n999), .C2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  AND4_X1   g576(.A1(new_n1001), .A2(new_n983), .A3(new_n994), .A4(new_n905), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(KEYINPUT43), .B2(new_n999), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(G397));
  AOI21_X1  g580(.A(G1384), .B1(new_n489), .B2(new_n493), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT112), .B(G40), .Z(new_n1009));
  NOR2_X1   g584(.A1(new_n473), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(KEYINPUT46), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT46), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  INV_X1    g590(.A(G2067), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n817), .B(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1011), .B1(new_n808), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  INV_X1    g595(.A(new_n736), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n734), .B(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1012), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n808), .B(G1996), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1011), .B1(new_n1025), .B2(new_n1017), .ZN(new_n1026));
  XOR2_X1   g601(.A(new_n1026), .B(KEYINPUT113), .Z(new_n1027));
  AND2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  OR3_X1    g603(.A1(G290), .A2(G1986), .A3(new_n1011), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1020), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n734), .A2(new_n1021), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT126), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G2067), .B2(new_n817), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1011), .B1(new_n1038), .B2(KEYINPUT127), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1010), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n706), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1010), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(KEYINPUT50), .B2(new_n1007), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1006), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1048), .A2(new_n1049), .B1(new_n1054), .B2(G2090), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT115), .B1(new_n1047), .B2(new_n706), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1044), .B(G8), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n690), .A2(new_n699), .ZN(new_n1058));
  OAI21_X1  g633(.A(G1981), .B1(new_n570), .B2(new_n574), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1058), .A2(KEYINPUT49), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1010), .B2(new_n1006), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n710), .A2(G1976), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1063), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n710), .B2(G1976), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1067), .B2(KEYINPUT52), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT116), .B(new_n1068), .C1(new_n1066), .C2(new_n1063), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1057), .A2(new_n1065), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1058), .B1(new_n1065), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1064), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1074), .A2(new_n1065), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1053), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1006), .A2(KEYINPUT118), .A3(new_n1052), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G2090), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1051), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1062), .B1(new_n1089), .B2(new_n1048), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1044), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1092), .A2(new_n1010), .A3(new_n1053), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1093), .A2(new_n796), .B1(new_n1047), .B2(new_n757), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1094), .A2(new_n1062), .A3(G286), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1083), .A2(new_n1091), .A3(new_n1057), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1095), .A2(KEYINPUT63), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1044), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND4_X1   g677(.A1(new_n1057), .A2(new_n1099), .A3(new_n1083), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1082), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G168), .A2(new_n1062), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT51), .B1(new_n1105), .B2(KEYINPUT123), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1106), .B(new_n1107), .C1(new_n1094), .C2(new_n1062), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1107), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1047), .A2(new_n757), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1051), .A2(new_n796), .A3(new_n1053), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1109), .B(G8), .C1(new_n1112), .C2(G286), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1105), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1108), .A2(new_n1113), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT124), .B(G1961), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1054), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1047), .B2(G2078), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1123), .B(new_n1125), .C1(new_n1047), .C2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1117), .A2(new_n1121), .A3(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n562), .A2(KEYINPUT119), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT57), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(new_n610), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1087), .B2(new_n1051), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(new_n792), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1047), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1139), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1087), .A2(new_n1051), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1141), .B(new_n1133), .C1(new_n1142), .C2(G1956), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1093), .A2(G1348), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1010), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n602), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1140), .B1(new_n1144), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1140), .A2(new_n1143), .A3(KEYINPUT61), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(KEYINPUT60), .C1(G1348), .C2(new_n1093), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1159), .A3(new_n602), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT58), .B(G1341), .Z(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1050), .B2(new_n1007), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1047), .B2(G1996), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(new_n552), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n552), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT122), .A3(new_n1169), .ZN(new_n1170));
  AND4_X1   g745(.A1(new_n1160), .A2(new_n1162), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1152), .B1(new_n1155), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1173));
  XNOR2_X1  g748(.A(G301), .B(KEYINPUT54), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1175));
  INV_X1    g750(.A(G40), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n473), .A2(new_n1176), .A3(new_n1126), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1173), .A2(new_n1178), .B1(new_n1127), .B2(new_n1174), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1116), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1130), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1083), .A2(new_n1091), .A3(new_n1057), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1104), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n722), .B(G1986), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1028), .B1(new_n1011), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1041), .B1(new_n1183), .B2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g761(.A1(G229), .A2(G227), .A3(new_n459), .A4(G401), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n906), .B2(new_n907), .ZN(new_n1189));
  NOR2_X1   g763(.A1(new_n1003), .A2(new_n1189), .ZN(G308));
  NAND3_X1  g764(.A1(new_n909), .A2(new_n905), .A3(new_n904), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1191), .B(new_n1188), .C1(new_n1192), .C2(new_n1002), .ZN(G225));
endmodule


