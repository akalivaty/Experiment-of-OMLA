//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT64), .A2(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT64), .A2(G134), .ZN(new_n190));
  OAI211_X1 g004(.A(new_n187), .B(new_n188), .C1(new_n189), .C2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(G134), .B2(new_n188), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n190), .ZN(new_n195));
  AOI21_X1  g009(.A(G131), .B1(new_n195), .B2(G137), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT65), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT65), .B1(new_n194), .B2(new_n196), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n197), .A2(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT0), .A4(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n203), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT0), .B(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G134), .ZN(new_n216));
  AOI21_X1  g030(.A(G137), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n192), .B1(new_n217), .B2(new_n187), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n216), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n201), .B1(new_n219), .B2(new_n188), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n224));
  OAI211_X1 g038(.A(G128), .B(new_n224), .C1(new_n208), .C2(new_n209), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n204), .B(new_n206), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n188), .A2(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n201), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n202), .A2(new_n213), .B1(new_n223), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G119), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G116), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G119), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(G113), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT2), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G113), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n238), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n240), .A2(new_n242), .A3(new_n238), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n237), .A2(KEYINPUT66), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G116), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(G119), .ZN(new_n249));
  INV_X1    g063(.A(new_n235), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n240), .A2(new_n242), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n240), .A2(new_n242), .A3(new_n238), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n233), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n259));
  INV_X1    g073(.A(new_n257), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n201), .B1(new_n194), .B2(new_n199), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n221), .B2(new_n222), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n212), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n232), .B1(new_n197), .B2(new_n198), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n259), .B(new_n260), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n202), .A2(new_n213), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(KEYINPUT69), .B(new_n232), .C1(new_n197), .C2(new_n198), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n267), .A2(new_n269), .A3(new_n257), .A4(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n264), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n260), .ZN(new_n276));
  NOR2_X1   g090(.A1(G237), .A2(G953), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G210), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n278), .B(KEYINPUT27), .Z(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G101), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n279), .B(new_n280), .Z(new_n281));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  INV_X1    g097(.A(new_n281), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n260), .B1(new_n233), .B2(KEYINPUT30), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n269), .A2(new_n270), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT30), .B1(new_n262), .B2(new_n212), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT70), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n202), .B2(new_n213), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n269), .A4(new_n270), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n285), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n271), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT73), .B(G902), .Z(new_n297));
  NOR2_X1   g111(.A1(new_n284), .A2(new_n283), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n260), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n274), .B1(new_n300), .B2(new_n271), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT72), .B(new_n274), .C1(new_n300), .C2(new_n271), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n296), .A2(new_n297), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G472), .ZN(new_n307));
  INV_X1    g121(.A(new_n285), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT69), .B1(new_n223), .B2(new_n232), .ZN(new_n309));
  INV_X1    g123(.A(new_n270), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n291), .B1(new_n311), .B2(new_n290), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT70), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT31), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n271), .A2(new_n281), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT31), .B1(new_n293), .B2(new_n316), .ZN(new_n319));
  INV_X1    g133(.A(new_n276), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n272), .B2(KEYINPUT28), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n318), .B(new_n319), .C1(new_n321), .C2(new_n281), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n323));
  NOR2_X1   g137(.A1(G472), .A2(G902), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n307), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT74), .B(G217), .Z(new_n328));
  INV_X1    g142(.A(new_n297), .ZN(new_n329));
  INV_X1    g143(.A(G234), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  INV_X1    g147(.A(G221), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n334), .A2(new_n330), .A3(G953), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n226), .A2(G119), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT23), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G119), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT23), .A2(G119), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT75), .B1(new_n346), .B2(G128), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(new_n226), .A3(KEYINPUT23), .A4(G119), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n337), .B1(new_n350), .B2(G110), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n345), .A2(new_n340), .ZN(new_n352));
  XOR2_X1   g166(.A(KEYINPUT24), .B(G110), .Z(new_n353));
  OR2_X1    g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g168(.A1(KEYINPUT76), .A2(new_n341), .B1(new_n226), .B2(G119), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n355), .A2(new_n339), .B1(new_n344), .B2(G128), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n347), .A2(new_n349), .ZN(new_n357));
  INV_X1    g171(.A(G110), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT77), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n354), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT16), .ZN(new_n361));
  INV_X1    g175(.A(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G125), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(G125), .ZN(new_n364));
  INV_X1    g178(.A(G125), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(G146), .B(new_n363), .C1(new_n367), .C2(new_n361), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n366), .A3(new_n203), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n363), .B1(new_n367), .B2(new_n361), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n203), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n368), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n350), .A2(G110), .B1(new_n352), .B2(new_n353), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n360), .A2(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n336), .B1(new_n375), .B2(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n360), .A2(new_n370), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n376), .B1(new_n383), .B2(new_n336), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT25), .B1(new_n384), .B2(new_n297), .ZN(new_n385));
  INV_X1    g199(.A(new_n336), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n381), .B2(new_n382), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n388));
  NOR4_X1   g202(.A1(new_n387), .A2(new_n388), .A3(new_n329), .A4(new_n376), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n332), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n332), .A2(G902), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n395));
  OAI21_X1  g209(.A(G214), .B1(G237), .B2(G902), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT83), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n212), .B2(G125), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n225), .A2(new_n227), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(G125), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n228), .A2(new_n398), .A3(new_n365), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT87), .B(G224), .Z(new_n404));
  INV_X1    g218(.A(G953), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n403), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n239), .B1(new_n235), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n251), .B2(new_n408), .ZN(new_n410));
  INV_X1    g224(.A(G101), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G104), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G107), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n412), .A3(KEYINPUT3), .A4(G104), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n414), .A2(KEYINPUT79), .A3(G107), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n412), .B2(G104), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n416), .B1(new_n422), .B2(new_n411), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n237), .A2(new_n252), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n422), .B2(new_n411), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n420), .B(new_n415), .C1(new_n413), .C2(KEYINPUT79), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(new_n429), .A3(G101), .A4(new_n418), .ZN(new_n430));
  OAI211_X1 g244(.A(G101), .B(new_n418), .C1(new_n419), .C2(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT80), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n427), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n426), .A3(G101), .A4(new_n418), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n245), .A2(new_n256), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n425), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n427), .A2(new_n430), .A3(new_n432), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n440), .A2(new_n256), .A3(new_n245), .A4(new_n434), .ZN(new_n441));
  INV_X1    g255(.A(new_n438), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n425), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n441), .B2(new_n425), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n445), .A2(new_n436), .A3(new_n447), .A4(new_n438), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n407), .B(new_n444), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT7), .B1(new_n406), .B2(KEYINPUT89), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(KEYINPUT89), .B2(new_n406), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n403), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT8), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n438), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n425), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n423), .B1(new_n410), .B2(new_n424), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT88), .B(KEYINPUT7), .Z(new_n459));
  NAND2_X1  g273(.A1(new_n406), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n401), .A2(new_n402), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n453), .A2(new_n443), .A3(new_n458), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G902), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n450), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G210), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n450), .A2(new_n466), .A3(new_n464), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n397), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G475), .ZN(new_n471));
  INV_X1    g285(.A(G237), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n405), .A3(G214), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT90), .A2(G143), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(KEYINPUT90), .A2(G143), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g291(.A1(KEYINPUT90), .A2(G143), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(G214), .A3(new_n277), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT18), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n201), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n367), .A2(G146), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n369), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n478), .A2(new_n474), .B1(new_n277), .B2(G214), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n473), .A2(new_n476), .ZN(new_n485));
  OAI21_X1  g299(.A(G131), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n481), .B(new_n483), .C1(new_n486), .C2(new_n480), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n484), .A2(new_n485), .A3(G131), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n201), .B1(new_n477), .B2(new_n479), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT17), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n372), .B(new_n368), .C1(new_n486), .C2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n487), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G113), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n414), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n495), .B(new_n487), .C1(new_n490), .C2(new_n492), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n471), .B1(new_n499), .B2(new_n463), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n488), .A2(new_n489), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT19), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT19), .B1(new_n364), .B2(new_n366), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n368), .B1(new_n504), .B2(G146), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n487), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n496), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n498), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT91), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n514));
  INV_X1    g328(.A(new_n510), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(KEYINPUT20), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n500), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G128), .B(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n195), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n205), .A2(G128), .ZN(new_n522));
  OAI21_X1  g336(.A(G134), .B1(new_n522), .B2(KEYINPUT13), .ZN(new_n523));
  AND2_X1   g337(.A1(KEYINPUT92), .A2(G122), .ZN(new_n524));
  NOR2_X1   g338(.A1(KEYINPUT92), .A2(G122), .ZN(new_n525));
  OAI21_X1  g339(.A(G116), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n246), .A2(new_n248), .A3(G122), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n526), .A2(new_n527), .A3(new_n412), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n412), .B1(new_n526), .B2(new_n527), .ZN(new_n529));
  OAI221_X1 g343(.A(new_n520), .B1(new_n521), .B2(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n226), .A2(G143), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n219), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n528), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n520), .A3(KEYINPUT93), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n527), .A2(KEYINPUT14), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT14), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n236), .A2(new_n541), .A3(G122), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n542), .A3(new_n526), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(G107), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n530), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT9), .B(G234), .Z(new_n546));
  NAND3_X1  g360(.A1(new_n328), .A2(new_n546), .A3(new_n405), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n530), .B(new_n549), .C1(new_n539), .C2(new_n544), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n329), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G478), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(KEYINPUT15), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n552), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n543), .A2(G107), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(new_n537), .A3(new_n538), .A4(new_n536), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n549), .B1(new_n558), .B2(new_n530), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n297), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n554), .A2(KEYINPUT15), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT95), .B(G952), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n329), .A2(G953), .A3(new_n565), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n555), .A2(new_n562), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n518), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n470), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n334), .B1(new_n546), .B2(new_n463), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G140), .ZN(new_n579));
  INV_X1    g393(.A(G227), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G953), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n579), .B(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n400), .A2(new_n423), .A3(KEYINPUT10), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n431), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n212), .B1(new_n426), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n440), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n400), .A2(new_n423), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n400), .A2(new_n423), .A3(KEYINPUT81), .A4(KEYINPUT10), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n585), .A2(new_n588), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n202), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n400), .A2(new_n423), .A3(KEYINPUT10), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n595), .A2(KEYINPUT81), .B1(new_n440), .B2(new_n587), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT10), .B1(new_n400), .B2(new_n423), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n584), .B2(new_n583), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n262), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n582), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n262), .B2(KEYINPUT82), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n400), .B(new_n423), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n202), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n598), .A3(new_n262), .ZN(new_n606));
  INV_X1    g420(.A(new_n582), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n603), .A2(new_n202), .A3(KEYINPUT82), .A4(new_n601), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n600), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G469), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n297), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n582), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n202), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n606), .A3(new_n607), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n611), .B1(new_n618), .B2(new_n463), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n578), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n395), .B1(new_n576), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n619), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n577), .B1(new_n622), .B2(new_n612), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT96), .A3(new_n575), .A4(new_n470), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n327), .A2(new_n394), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND2_X1  g440(.A1(new_n322), .A2(new_n297), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(G472), .B1(new_n324), .B2(new_n322), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n620), .A2(new_n393), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  OAI22_X1  g447(.A1(new_n556), .A2(new_n559), .B1(KEYINPUT97), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n551), .A2(new_n552), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n297), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G478), .ZN(new_n639));
  AOI211_X1 g453(.A(G478), .B(new_n329), .C1(new_n551), .C2(new_n552), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n632), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI211_X1 g456(.A(KEYINPUT98), .B(new_n640), .C1(new_n638), .C2(G478), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n642), .A2(new_n643), .A3(new_n518), .ZN(new_n644));
  INV_X1    g458(.A(new_n396), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n468), .B2(new_n469), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n644), .A2(KEYINPUT99), .A3(new_n572), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n639), .A2(new_n641), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n514), .A2(new_n517), .ZN(new_n651));
  INV_X1    g465(.A(new_n500), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n639), .A2(new_n632), .A3(new_n641), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n450), .A2(new_n466), .A3(new_n464), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n466), .B1(new_n450), .B2(new_n464), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n572), .B(new_n396), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n648), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n647), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n631), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  XNOR2_X1  g477(.A(new_n513), .B(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n555), .A2(new_n562), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n666), .A3(new_n652), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n631), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NOR2_X1   g485(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n379), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n391), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n390), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n621), .A2(new_n624), .A3(new_n628), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT100), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G12));
  OAI21_X1  g493(.A(new_n566), .B1(new_n568), .B2(G900), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n667), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n390), .A2(new_n674), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n396), .B1(new_n656), .B2(new_n657), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n683), .A2(new_n620), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n327), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XNOR2_X1  g501(.A(new_n680), .B(KEYINPUT39), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n623), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT40), .Z(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n665), .B1(new_n651), .B2(new_n652), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n396), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n691), .B1(new_n694), .B2(new_n683), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n693), .A2(new_n675), .A3(KEYINPUT101), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n656), .A2(new_n657), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n293), .A2(new_n294), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n284), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n300), .A2(new_n271), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n463), .B1(new_n702), .B2(new_n281), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n325), .B2(new_n326), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n690), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR4_X1   g521(.A1(new_n642), .A2(new_n643), .A3(new_n518), .A4(new_n681), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n327), .A2(new_n685), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AND4_X1   g524(.A1(new_n606), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n607), .B1(new_n616), .B2(new_n606), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n297), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(KEYINPUT102), .A2(G469), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n610), .A2(new_n297), .A3(new_n714), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n578), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT103), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n660), .A2(new_n327), .A3(new_n394), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT104), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  NAND4_X1  g537(.A1(new_n327), .A2(new_n668), .A3(new_n394), .A4(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  OAI21_X1  g539(.A(KEYINPUT105), .B1(new_n684), .B2(new_n718), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n714), .B1(new_n610), .B2(new_n297), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n329), .B(new_n715), .C1(new_n600), .C2(new_n609), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n577), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n646), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n675), .A2(new_n575), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n327), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n327), .A2(KEYINPUT106), .A3(new_n732), .A4(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  NAND2_X1  g553(.A1(new_n646), .A2(new_n692), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n571), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT72), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n702), .A2(new_n742), .A3(KEYINPUT28), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n301), .B2(new_n302), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n319), .B(new_n318), .C1(new_n744), .C2(new_n281), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n627), .A2(G472), .B1(new_n324), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n719), .A2(new_n741), .A3(new_n746), .A4(new_n394), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NAND4_X1  g562(.A1(new_n732), .A2(new_n675), .A3(new_n708), .A4(new_n746), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NOR3_X1   g564(.A1(new_n656), .A2(new_n657), .A3(new_n645), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n615), .B2(new_n617), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n617), .A2(new_n753), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n611), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n611), .A2(new_n463), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n612), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n578), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n327), .A2(new_n394), .A3(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  INV_X1    g579(.A(new_n708), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n763), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n763), .B(KEYINPUT42), .C1(new_n762), .C2(new_n766), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND4_X1  g585(.A1(new_n327), .A2(new_n394), .A3(new_n682), .A4(new_n761), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NOR2_X1   g587(.A1(new_n628), .A2(new_n683), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n642), .A2(new_n643), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n653), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(KEYINPUT110), .B2(KEYINPUT43), .ZN(new_n778));
  AND2_X1   g592(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n779));
  NOR2_X1   g593(.A1(KEYINPUT110), .A2(KEYINPUT43), .ZN(new_n780));
  OAI22_X1  g594(.A1(new_n776), .A2(new_n653), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n778), .A2(KEYINPUT111), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n778), .B2(new_n781), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n774), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n752), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n688), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n754), .A2(new_n788), .A3(new_n755), .ZN(new_n789));
  INV_X1    g603(.A(new_n618), .ZN(new_n790));
  OAI21_X1  g604(.A(G469), .B1(new_n790), .B2(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n758), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT109), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n613), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n577), .B(new_n787), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n786), .B(new_n797), .C1(new_n785), .C2(new_n784), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  NOR4_X1   g613(.A1(new_n327), .A2(new_n766), .A3(new_n394), .A4(new_n752), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n796), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(KEYINPUT47), .A3(new_n578), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT47), .B1(new_n801), .B2(new_n578), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  NOR2_X1   g619(.A1(new_n577), .A2(new_n397), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n777), .A2(new_n394), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n705), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n716), .A2(new_n717), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT49), .Z(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n698), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n623), .A2(new_n646), .A3(new_n675), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n318), .A2(new_n319), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n321), .A2(new_n281), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n324), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT32), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n813), .B1(new_n819), .B2(new_n307), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n627), .A2(G472), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n745), .A2(new_n324), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n821), .A2(new_n708), .A3(new_n675), .A4(new_n822), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n820), .A2(new_n682), .B1(new_n823), .B2(new_n732), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n390), .A2(new_n674), .A3(new_n680), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n740), .A2(new_n760), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n820), .A2(new_n708), .B1(new_n705), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n705), .A2(new_n826), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n686), .A2(new_n709), .A3(new_n749), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT114), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(new_n829), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n761), .A2(new_n746), .A3(new_n675), .A4(new_n708), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n652), .A2(new_n664), .A3(new_n665), .A4(new_n680), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n623), .A2(new_n837), .A3(new_n675), .A4(new_n751), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n327), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n772), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n768), .A2(new_n769), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n720), .A2(new_n724), .A3(new_n747), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n738), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n470), .A2(new_n572), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n518), .A2(new_n666), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n655), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n628), .A3(new_n629), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n625), .A2(new_n676), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT112), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n625), .A2(new_n676), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n844), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n812), .B1(new_n835), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n828), .B1(new_n824), .B2(new_n827), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n831), .A2(KEYINPUT114), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n686), .A2(new_n749), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT113), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n812), .B1(new_n850), .B2(new_n852), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n841), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n842), .A2(new_n867), .A3(new_n738), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n867), .B1(new_n842), .B2(new_n738), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n866), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g686(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n855), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n835), .A2(new_n854), .A3(KEYINPUT115), .A4(new_n812), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n829), .A2(new_n832), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n856), .A2(new_n876), .B1(new_n861), .B2(new_n862), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n812), .B1(new_n877), .B2(new_n854), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT115), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n850), .A2(new_n852), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n768), .A2(new_n840), .A3(new_n769), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n843), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n829), .A2(new_n832), .A3(KEYINPUT52), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n859), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT53), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n875), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n874), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n752), .A2(new_n393), .A3(new_n566), .A4(new_n718), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n808), .A2(new_n644), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n564), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n566), .B1(new_n778), .B2(new_n781), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n893), .A2(new_n394), .A3(new_n746), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n894), .B2(new_n732), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n752), .A2(new_n718), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT48), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n327), .A2(new_n394), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n898), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n895), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n898), .A2(new_n675), .A3(new_n746), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n698), .A2(new_n645), .A3(new_n729), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n894), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT50), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n894), .A2(KEYINPUT50), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n808), .A2(new_n518), .A3(new_n776), .A4(new_n890), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n802), .A2(new_n803), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n578), .B2(new_n809), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n751), .A3(new_n894), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n905), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n906), .A2(new_n912), .A3(KEYINPUT119), .A4(new_n913), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n924), .B2(KEYINPUT51), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n889), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n811), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n405), .A2(G952), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n407), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n883), .B2(new_n885), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(new_n841), .A3(new_n865), .A4(new_n868), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n935), .A2(new_n877), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n329), .B(new_n467), .C1(new_n933), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n329), .B1(new_n933), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT120), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n942), .B(new_n329), .C1(new_n933), .C2(new_n936), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n467), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n932), .A2(new_n938), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n929), .B(new_n939), .C1(new_n944), .C2(new_n945), .ZN(G51));
  INV_X1    g760(.A(new_n873), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n933), .A2(new_n936), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n873), .B1(new_n855), .B2(new_n872), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n757), .B(KEYINPUT57), .Z(new_n951));
  OAI21_X1  g765(.A(new_n610), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n791), .A2(new_n789), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n941), .A2(new_n953), .A3(new_n943), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n929), .B1(new_n952), .B2(new_n954), .ZN(G54));
  NAND2_X1  g769(.A1(KEYINPUT58), .A2(G475), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT121), .Z(new_n957));
  NAND3_X1  g771(.A1(new_n941), .A2(new_n943), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n512), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n511), .B1(new_n507), .B2(new_n498), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n958), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n929), .ZN(G60));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  INV_X1    g780(.A(new_n929), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n634), .A2(new_n637), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT59), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n966), .B(new_n967), .C1(new_n950), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n947), .B1(new_n933), .B2(new_n936), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(new_n874), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT122), .B1(new_n974), .B2(new_n929), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n968), .B1(new_n889), .B2(new_n970), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G63));
  XOR2_X1   g792(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n979));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n855), .B2(new_n872), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT124), .B(new_n967), .C1(new_n982), .C2(new_n384), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n673), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n981), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n933), .B2(new_n936), .ZN(new_n987));
  INV_X1    g801(.A(new_n384), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT124), .B1(new_n989), .B2(new_n967), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n979), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n929), .B1(new_n987), .B2(new_n988), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n984), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT125), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n992), .A2(new_n995), .A3(KEYINPUT61), .A4(new_n984), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(G66));
  INV_X1    g811(.A(new_n404), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n998), .B2(new_n570), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n881), .A2(new_n843), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n930), .B1(G898), .B2(new_n405), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G69));
  OAI22_X1  g817(.A1(new_n312), .A2(new_n313), .B1(KEYINPUT30), .B2(new_n233), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(new_n504), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(G900), .B(G953), .C1(new_n1006), .C2(G227), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(G227), .B2(new_n1006), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n860), .A2(KEYINPUT113), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n860), .A2(KEYINPUT113), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n1009), .A2(new_n1010), .B1(new_n820), .B2(new_n708), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n706), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n804), .A2(new_n798), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n655), .A2(new_n846), .ZN(new_n1018));
  NOR4_X1   g832(.A1(new_n900), .A2(new_n689), .A3(new_n752), .A4(new_n1018), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n1005), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n797), .A2(new_n901), .A3(new_n646), .A4(new_n692), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1023), .A2(new_n770), .A3(new_n772), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1011), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1017), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(G953), .B1(new_n1026), .B2(new_n1006), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1008), .B1(new_n1022), .B2(new_n1027), .ZN(G72));
  INV_X1    g842(.A(new_n701), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1015), .A2(new_n1000), .A3(new_n1020), .ZN(new_n1030));
  XOR2_X1   g844(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n1031));
  NAND2_X1  g845(.A1(G472), .A2(G902), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n700), .A2(new_n284), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1029), .A2(new_n1035), .A3(new_n1033), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n887), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1026), .A2(new_n1000), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1035), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  NOR4_X1   g853(.A1(new_n1034), .A2(new_n1037), .A3(new_n1039), .A4(new_n929), .ZN(G57));
endmodule


