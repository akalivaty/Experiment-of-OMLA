//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT78), .A2(G104), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT78), .A2(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(G104), .A2(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G101), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT80), .B(G101), .Z(new_n195));
  OAI22_X1  g009(.A1(new_n188), .A2(new_n189), .B1(KEYINPUT3), .B2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT3), .A2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n187), .A3(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n190), .A2(KEYINPUT81), .A3(G101), .A4(new_n191), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT83), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(KEYINPUT83), .A3(new_n200), .A4(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .A4(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(KEYINPUT67), .A3(new_n211), .A4(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT68), .A2(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT68), .A2(G128), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n208), .A2(new_n210), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT10), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n200), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n196), .A2(new_n197), .A3(new_n199), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n229), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT0), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n222), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n215), .B1(new_n236), .B2(new_n237), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n206), .A2(new_n226), .B1(new_n234), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n194), .A2(new_n200), .A3(new_n201), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n218), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n222), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n217), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT82), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n214), .A2(new_n216), .B1(new_n222), .B2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n202), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n243), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  OAI211_X1 g068(.A(G134), .B(new_n253), .C1(new_n254), .C2(KEYINPUT65), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(KEYINPUT11), .C1(new_n257), .C2(G137), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  AOI22_X1  g074(.A1(KEYINPUT65), .A2(new_n254), .B1(new_n257), .B2(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n242), .A2(new_n252), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n242), .A2(new_n252), .A3(KEYINPUT84), .A4(new_n265), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n194), .A2(new_n201), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(KEYINPUT82), .A3(new_n247), .A4(new_n200), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n250), .B1(new_n202), .B2(new_n249), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT10), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n234), .A2(new_n241), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n225), .B1(new_n204), .B2(new_n205), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n277), .A2(new_n265), .ZN(new_n278));
  XNOR2_X1  g092(.A(G110), .B(G140), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT77), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G227), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n270), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  OAI22_X1  g098(.A1(new_n248), .A2(new_n251), .B1(new_n224), .B2(new_n244), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(KEYINPUT12), .C1(new_n264), .C2(new_n263), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n214), .A2(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n272), .A2(new_n273), .B1(new_n288), .B2(new_n202), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n289), .B2(new_n265), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n268), .A2(new_n269), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n284), .B(G469), .C1(new_n283), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(G469), .A2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n290), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n270), .A2(new_n283), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n283), .B1(new_n270), .B2(new_n278), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n295), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT84), .B1(new_n277), .B2(new_n265), .ZN(new_n303));
  INV_X1    g117(.A(new_n269), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n283), .B(new_n297), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n277), .A2(new_n265), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n268), .B2(new_n269), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n307), .B2(new_n283), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT85), .A3(new_n295), .A4(new_n296), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n294), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n239), .B2(new_n240), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n224), .B2(new_n311), .ZN(new_n313));
  INV_X1    g127(.A(G224), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT7), .B1(new_n314), .B2(G953), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT88), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n314), .A2(G953), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n313), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G116), .B(G119), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT2), .B(G113), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G119), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT5), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n324), .A2(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G113), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n322), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n202), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G122), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT8), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n319), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n320), .A2(new_n321), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n332), .B(new_n334), .C1(new_n202), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n281), .A2(G224), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n241), .A2(G125), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n288), .B2(G125), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT7), .B(new_n342), .C1(new_n344), .C2(KEYINPUT88), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n318), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n319), .B(new_n321), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n206), .A2(new_n331), .B1(new_n234), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n333), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n318), .A2(new_n345), .A3(new_n341), .A4(KEYINPUT89), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n296), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n351), .A2(new_n333), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT6), .A3(new_n352), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n313), .B(new_n317), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n333), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n354), .A2(KEYINPUT90), .A3(new_n296), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n357), .A2(new_n367), .A3(new_n364), .A4(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT9), .B(G234), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n310), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n281), .A2(G221), .A3(G234), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT22), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(G137), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT75), .ZN(new_n382));
  XOR2_X1   g196(.A(G125), .B(G140), .Z(new_n383));
  OAI21_X1  g197(.A(KEYINPUT73), .B1(new_n383), .B2(G146), .ZN(new_n384));
  XNOR2_X1  g198(.A(G125), .B(G140), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n207), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n384), .A2(new_n387), .B1(new_n389), .B2(G146), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n323), .B1(new_n219), .B2(new_n220), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n237), .A2(G119), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(KEYINPUT23), .A3(new_n394), .ZN(new_n395));
  OR3_X1    g209(.A1(new_n323), .A2(KEYINPUT23), .A3(G128), .ZN(new_n396));
  AOI21_X1  g210(.A(G110), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT24), .B(G110), .Z(new_n398));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n392), .A2(new_n399), .A3(new_n394), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT72), .B1(new_n391), .B2(new_n393), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n390), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n388), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n383), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n207), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n389), .A2(G146), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n395), .A2(G110), .A3(new_n396), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n401), .A3(new_n398), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT74), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n403), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n403), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n382), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n403), .A2(new_n412), .A3(new_n381), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(new_n296), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT25), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n416), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(G234), .B2(new_n296), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(KEYINPUT76), .A3(new_n424), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n416), .A2(new_n417), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n424), .A2(G902), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n434));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n253), .A2(G134), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n257), .A2(G137), .ZN(new_n437));
  OAI21_X1  g251(.A(G131), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n262), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n435), .B1(new_n262), .B2(new_n438), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n288), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n241), .B1(new_n263), .B2(new_n264), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n434), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n224), .A2(new_n262), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n442), .A3(KEYINPUT30), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n350), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n442), .A3(new_n349), .ZN(new_n448));
  NOR2_X1   g262(.A1(G237), .A2(G953), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G210), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT27), .Z(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT26), .ZN(new_n452));
  INV_X1    g266(.A(G101), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n448), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT69), .B1(new_n455), .B2(KEYINPUT31), .ZN(new_n456));
  INV_X1    g270(.A(new_n448), .ZN(new_n457));
  INV_X1    g271(.A(new_n434), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n262), .A2(new_n438), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n262), .A2(new_n435), .A3(new_n438), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n224), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n442), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n457), .B1(new_n465), .B2(new_n350), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT31), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n454), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n456), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n457), .A2(KEYINPUT28), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n448), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n350), .B1(new_n441), .B2(new_n443), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n454), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n455), .A2(KEYINPUT31), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G472), .A2(G902), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT32), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n481));
  INV_X1    g295(.A(new_n479), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n481), .B(new_n482), .C1(new_n470), .C2(new_n477), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT70), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n466), .B2(new_n454), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT29), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n447), .A2(new_n448), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(KEYINPUT70), .A3(new_n476), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n487), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n288), .A2(new_n459), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n350), .B1(new_n443), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n448), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n445), .A2(KEYINPUT71), .A3(new_n442), .A4(new_n349), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(KEYINPUT28), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n497), .A2(KEYINPUT29), .A3(new_n454), .A4(new_n473), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(new_n296), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G472), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n433), .B1(new_n484), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n375), .A2(new_n423), .A3(G953), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n219), .A2(new_n220), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G143), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n505), .A2(KEYINPUT13), .B1(G128), .B2(new_n209), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n209), .A2(KEYINPUT13), .A3(G128), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT96), .Z(new_n508));
  OAI21_X1  g322(.A(G134), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n510), .A2(KEYINPUT95), .A3(G116), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT95), .B1(new_n510), .B2(G116), .ZN(new_n512));
  OAI22_X1  g326(.A1(new_n511), .A2(new_n512), .B1(G116), .B2(new_n510), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(G107), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n209), .A2(G128), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n505), .A2(new_n257), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n509), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT97), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n505), .A2(new_n515), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G134), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n516), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(new_n511), .B2(new_n512), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n513), .A2(new_n525), .A3(G107), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n187), .A2(KEYINPUT14), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n503), .B1(new_n521), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  INV_X1    g345(.A(new_n503), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n531), .B(new_n532), .C1(new_n519), .C2(new_n520), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n296), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G478), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI221_X1 g351(.A(new_n296), .B1(KEYINPUT15), .B2(new_n535), .C1(new_n530), .C2(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n409), .ZN(new_n540));
  INV_X1    g354(.A(G237), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n281), .A3(G214), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n209), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n449), .B(G214), .C1(KEYINPUT91), .C2(G143), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT17), .A3(G131), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(G131), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n540), .B(new_n547), .C1(KEYINPUT17), .C2(new_n548), .ZN(new_n549));
  XOR2_X1   g363(.A(G113), .B(G122), .Z(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G104), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n546), .A2(KEYINPUT92), .A3(KEYINPUT18), .A4(G131), .ZN(new_n552));
  AND3_X1   g366(.A1(KEYINPUT92), .A2(KEYINPUT18), .A3(G131), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n384), .A2(new_n387), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n385), .A2(new_n207), .ZN(new_n555));
  OAI221_X1 g369(.A(new_n552), .B1(new_n546), .B2(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n549), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n551), .B1(new_n549), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n296), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT94), .B(new_n296), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(G475), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G475), .ZN(new_n564));
  OR3_X1    g378(.A1(new_n383), .A2(KEYINPUT93), .A3(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT93), .B1(new_n383), .B2(KEYINPUT19), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n548), .B(new_n408), .C1(new_n568), .C2(G146), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n551), .B1(new_n556), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n564), .B(new_n296), .C1(new_n557), .C2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n563), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(G234), .A2(G237), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(G952), .A3(new_n281), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT21), .B(G898), .Z(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n576), .A2(G902), .A3(G953), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n539), .A2(new_n575), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n378), .A2(new_n502), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT98), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n195), .ZN(G3));
  NOR3_X1   g401(.A1(new_n310), .A2(new_n433), .A3(new_n377), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n470), .B2(new_n477), .ZN(new_n589));
  INV_X1    g403(.A(G472), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT99), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT100), .Z(new_n594));
  NAND3_X1  g408(.A1(new_n369), .A2(KEYINPUT101), .A3(new_n370), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n521), .A2(new_n529), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n532), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n521), .A2(new_n529), .A3(new_n503), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(KEYINPUT33), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n530), .B2(new_n533), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n535), .A2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n534), .A2(new_n535), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n583), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n605), .A2(new_n575), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n366), .A2(new_n608), .A3(new_n368), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n372), .A2(new_n595), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n594), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  AND3_X1   g428(.A1(new_n595), .A2(new_n372), .A3(new_n609), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n575), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n583), .B(KEYINPUT102), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n539), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n594), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT35), .B(G107), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  INV_X1    g437(.A(new_n592), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT76), .B1(new_n422), .B2(new_n424), .ZN(new_n625));
  INV_X1    g439(.A(new_n424), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n426), .B(new_n626), .C1(new_n420), .C2(new_n421), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n414), .A2(new_n415), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n382), .A2(KEYINPUT36), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n628), .B(new_n629), .Z(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(new_n431), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n625), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n378), .A2(new_n584), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT103), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT37), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(G110), .Z(G12));
  NAND2_X1  g451(.A1(new_n302), .A2(new_n309), .ZN(new_n638));
  INV_X1    g452(.A(new_n294), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n377), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n632), .B1(new_n484), .B2(new_n501), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n617), .A2(new_n539), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n577), .B(KEYINPUT104), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n581), .A2(G900), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n640), .A2(new_n615), .A3(new_n641), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  AND2_X1   g463(.A1(new_n369), .A2(new_n370), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT38), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n539), .A2(new_n575), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n632), .A2(new_n372), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT105), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n455), .A2(KEYINPUT31), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n475), .A2(new_n476), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n456), .B2(new_n469), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n481), .B1(new_n661), .B2(new_n482), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n478), .A2(KEYINPUT32), .A3(new_n479), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n495), .A2(new_n496), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n296), .B1(new_n664), .B2(new_n454), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n466), .A2(new_n476), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n662), .A2(new_n663), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n645), .B(KEYINPUT39), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n640), .B2(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n640), .A2(KEYINPUT40), .A3(new_n670), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n657), .B(new_n669), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND3_X1  g488(.A1(new_n605), .A2(new_n575), .A3(new_n645), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n640), .A2(new_n615), .A3(new_n641), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI21_X1  g492(.A(new_n295), .B1(new_n308), .B2(new_n296), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n377), .B(new_n679), .C1(new_n302), .C2(new_n309), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n610), .A2(new_n680), .A3(new_n502), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  AND2_X1   g497(.A1(new_n574), .A2(new_n573), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n539), .A2(new_n684), .A3(new_n563), .A4(new_n619), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n372), .A2(new_n595), .A3(new_n609), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n680), .A3(new_n502), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND3_X1  g502(.A1(new_n662), .A2(new_n663), .A3(new_n501), .ZN(new_n689));
  INV_X1    g503(.A(new_n631), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n427), .A2(new_n690), .A3(new_n428), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n689), .A2(new_n584), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n680), .A3(new_n615), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  NAND4_X1  g508(.A1(new_n595), .A2(new_n372), .A3(new_n609), .A4(new_n652), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n497), .A2(new_n473), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n497), .A2(KEYINPUT106), .A3(new_n473), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n476), .A3(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(new_n470), .A3(new_n658), .ZN(new_n702));
  OAI22_X1  g516(.A1(new_n702), .A2(new_n482), .B1(new_n589), .B2(new_n590), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n433), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n696), .A2(new_n680), .A3(new_n619), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR3_X1   g520(.A1(new_n632), .A2(new_n703), .A3(new_n675), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n680), .A2(new_n707), .A3(new_n615), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT108), .B1(new_n711), .B2(new_n689), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n502), .A2(KEYINPUT108), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n293), .B(KEYINPUT107), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n638), .A2(new_n292), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n372), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n371), .A2(new_n377), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n676), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n502), .A3(new_n719), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n710), .B1(new_n724), .B2(new_n675), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n689), .A2(new_n711), .A3(KEYINPUT108), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT42), .B1(new_n726), .B2(new_n712), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT109), .B1(new_n727), .B2(new_n720), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND4_X1  g544(.A1(new_n717), .A2(new_n502), .A3(new_n647), .A4(new_n719), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  AND3_X1   g546(.A1(new_n270), .A2(new_n278), .A3(new_n283), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n283), .B1(new_n270), .B2(new_n297), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT45), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n733), .B2(new_n734), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(G469), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n716), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n716), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n638), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n376), .A3(new_n670), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  INV_X1    g562(.A(new_n605), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n748), .B1(new_n749), .B2(new_n575), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n617), .A2(KEYINPUT43), .A3(new_n605), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n624), .A2(new_n752), .A3(new_n691), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n650), .A2(new_n372), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n753), .B2(new_n754), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n376), .A4(new_n670), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n747), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NAND2_X1  g574(.A1(new_n744), .A2(new_n376), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n711), .A2(new_n689), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n744), .A2(new_n764), .A3(new_n376), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n756), .A2(new_n675), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n763), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  INV_X1    g582(.A(new_n679), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n638), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n756), .A3(new_n377), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n643), .B1(new_n750), .B2(new_n751), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n726), .A2(new_n712), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT48), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n680), .A2(new_n704), .A3(new_n772), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n616), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT118), .Z(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(KEYINPUT48), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n281), .A2(G952), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n669), .A2(new_n433), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n771), .A2(new_n578), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n605), .A2(new_n575), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n777), .A2(new_n780), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n632), .A2(new_n703), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n773), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT116), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n784), .A2(new_n617), .A3(new_n749), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n762), .A2(new_n765), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n376), .B2(new_n770), .ZN(new_n796));
  INV_X1    g610(.A(new_n756), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n704), .A3(new_n797), .A4(new_n772), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  INV_X1    g614(.A(new_n651), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n778), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n802), .B2(new_n718), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT50), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n804), .A2(KEYINPUT51), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n787), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n804), .A2(new_n809), .A3(new_n805), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n794), .A2(new_n798), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n804), .B2(new_n805), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n648), .A2(new_n677), .A3(new_n708), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n696), .A2(new_n376), .A3(new_n669), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n717), .A2(new_n632), .A3(new_n645), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n689), .A2(new_n691), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n310), .A3(new_n377), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n821), .B(new_n615), .C1(new_n647), .C2(new_n676), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n695), .A2(new_n377), .A3(new_n668), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n302), .A2(new_n309), .B1(G469), .B2(new_n735), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n691), .B1(new_n824), .B2(new_n716), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n645), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n708), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n819), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n785), .B1(new_n620), .B2(KEYINPUT111), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n830), .B(new_n718), .C1(new_n369), .C2(new_n370), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n831), .B2(new_n642), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n373), .B2(new_n618), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n588), .A2(new_n832), .A3(new_n592), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n585), .A3(new_n634), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n705), .A2(new_n681), .A3(new_n687), .A4(new_n693), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n539), .A2(new_n575), .A3(new_n646), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n640), .A2(new_n797), .A3(new_n641), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n717), .A2(new_n676), .A3(new_n788), .A4(new_n719), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n731), .A3(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n835), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n828), .A2(new_n841), .A3(new_n729), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT54), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n843), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  INV_X1    g663(.A(new_n840), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(KEYINPUT53), .C1(new_n836), .C2(KEYINPUT113), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n835), .B1(KEYINPUT113), .B2(new_n836), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n729), .A3(new_n828), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n843), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n848), .A2(new_n849), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n807), .A2(new_n813), .A3(new_n845), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(G952), .B2(G953), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n770), .B(KEYINPUT49), .Z(new_n859));
  NOR4_X1   g673(.A1(new_n749), .A2(new_n575), .A3(new_n377), .A4(new_n718), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n651), .A3(new_n783), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n861), .ZN(G75));
  NAND3_X1  g676(.A1(new_n848), .A2(new_n854), .A3(new_n855), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n359), .A2(new_n363), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n362), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT55), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n281), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G51));
  XOR2_X1   g686(.A(new_n716), .B(KEYINPUT57), .Z(new_n873));
  AND3_X1   g687(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n843), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT112), .B1(new_n842), .B2(new_n843), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n849), .B1(new_n876), .B2(new_n854), .ZN(new_n877));
  INV_X1    g691(.A(new_n856), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n308), .B(KEYINPUT119), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n739), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n863), .A2(G902), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n871), .B1(new_n881), .B2(new_n883), .ZN(G54));
  NAND4_X1  g698(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n557), .A2(new_n570), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n887), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n888), .A2(new_n889), .A3(new_n871), .ZN(G60));
  INV_X1    g704(.A(new_n871), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT59), .Z(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n845), .B2(new_n856), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n599), .A2(new_n601), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n877), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n897), .B2(new_n856), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n895), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT120), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n863), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n429), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n863), .A2(new_n630), .A3(new_n902), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n871), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n430), .B1(new_n863), .B2(new_n902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n891), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n907), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n580), .B2(new_n314), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n835), .A2(new_n836), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n866), .B1(G898), .B2(new_n281), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  NAND4_X1  g736(.A1(new_n759), .A2(new_n767), .A3(new_n729), .A4(new_n731), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n747), .A2(new_n696), .A3(new_n775), .A4(new_n758), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n815), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n822), .A2(KEYINPUT122), .A3(new_n708), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n281), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n281), .A2(G900), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n465), .B(new_n568), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n640), .A2(new_n670), .ZN(new_n934));
  INV_X1    g748(.A(new_n642), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n502), .B1(new_n935), .B2(new_n785), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n936), .A3(new_n756), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n673), .A2(new_n926), .A3(new_n927), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n673), .A2(new_n927), .A3(new_n926), .A4(KEYINPUT62), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n759), .A2(new_n767), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n932), .A2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n932), .A2(KEYINPUT124), .ZN(new_n947));
  NAND2_X1  g761(.A1(G227), .A2(G900), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(G953), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n946), .B(new_n949), .ZN(G72));
  NOR3_X1   g764(.A1(new_n923), .A2(new_n928), .A3(new_n918), .ZN(new_n951));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n466), .B(new_n476), .C1(new_n951), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n891), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n955), .B2(new_n891), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n942), .A2(new_n919), .A3(new_n943), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n953), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(KEYINPUT125), .A3(new_n953), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n963), .A2(new_n666), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n486), .A2(new_n455), .A3(new_n490), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n844), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n959), .A2(new_n965), .A3(new_n969), .ZN(G57));
endmodule


