//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n461), .B2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n466), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n460), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(new_n475), .A3(G125), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(KEYINPUT67), .A3(G125), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n473), .B1(G2105), .B2(new_n482), .ZN(G160));
  AOI21_X1  g058(.A(new_n466), .B1(new_n462), .B2(new_n464), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n462), .B2(new_n464), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G136), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n466), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n466), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n465), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n474), .A2(new_n475), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n466), .C1(new_n499), .C2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n494), .B(new_n498), .C1(new_n502), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XOR2_X1   g091(.A(new_n516), .B(KEYINPUT74), .Z(new_n517));
  OAI21_X1  g092(.A(new_n511), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n514), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  INV_X1    g103(.A(new_n526), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n510), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G543), .ZN(new_n531));
  OAI221_X1 g106(.A(new_n518), .B1(new_n519), .B2(new_n527), .C1(new_n528), .C2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  INV_X1    g108(.A(new_n531), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  INV_X1    g110(.A(new_n527), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  INV_X1    g112(.A(new_n514), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n521), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n539), .A2(G63), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n535), .A2(new_n537), .A3(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n534), .A2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n536), .A2(G90), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n510), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n510), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n530), .A2(G43), .A3(G543), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n527), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  OAI211_X1 g137(.A(G53), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n530), .A2(new_n565), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g142(.A(G91), .B(new_n514), .C1(new_n525), .C2(new_n526), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n530), .A2(new_n570), .A3(G91), .A4(new_n514), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n538), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n567), .A2(new_n572), .A3(new_n576), .ZN(G299));
  NAND3_X1  g152(.A1(new_n530), .A2(G87), .A3(new_n514), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n530), .A2(G49), .A3(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n582), .B(G651), .C1(new_n514), .C2(G74), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n578), .A2(new_n579), .A3(new_n581), .A4(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n530), .A2(G86), .A3(new_n514), .ZN(new_n585));
  OAI211_X1 g160(.A(G48), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n512), .B2(new_n513), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n511), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT77), .ZN(G305));
  NAND2_X1  g167(.A1(new_n536), .A2(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n534), .A2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n510), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g173(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n510), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  OAI211_X1 g176(.A(G54), .B(G543), .C1(new_n525), .C2(new_n526), .ZN(new_n602));
  OR2_X1    g177(.A1(KEYINPUT79), .A2(G66), .ZN(new_n603));
  NAND2_X1  g178(.A1(KEYINPUT79), .A2(G66), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(new_n514), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n602), .B1(new_n606), .B2(new_n521), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n527), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .A4(new_n514), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n601), .B1(G868), .B2(new_n612), .ZN(G284));
  OAI21_X1  g188(.A(new_n601), .B1(G868), .B2(new_n612), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n556), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n610), .A2(new_n611), .ZN(new_n623));
  INV_X1    g198(.A(new_n607), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n625), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n622), .B1(new_n626), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n471), .A2(new_n479), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(G2100), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n630), .ZN(new_n634));
  OR3_X1    g209(.A1(new_n634), .A2(new_n632), .A3(G2100), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n632), .B2(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n485), .A2(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n490), .B2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n636), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n654), .A2(new_n658), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT83), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n666), .B(KEYINPUT17), .Z(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n663), .A3(new_n667), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n663), .A3(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1971), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(G6), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n591), .B(KEYINPUT77), .Z(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n698), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT32), .B(G1981), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  MUX2_X1   g282(.A(G23), .B(G288), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n701), .A2(new_n706), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G25), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n490), .A2(G131), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT85), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n485), .A2(G119), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n715), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n723), .A2(new_n725), .ZN(new_n727));
  INV_X1    g302(.A(G24), .ZN(new_n728));
  OR3_X1    g303(.A1(new_n728), .A2(KEYINPUT87), .A3(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT87), .B1(new_n728), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G290), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n698), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1986), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n726), .A2(new_n727), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n712), .A2(new_n713), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT36), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n714), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n485), .A2(G129), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT92), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n490), .A2(G141), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n471), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n737), .B1(new_n746), .B2(new_n714), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT27), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G1996), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n698), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n698), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G1966), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n698), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n698), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1961), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n714), .B1(new_n756), .B2(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G160), .B2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2084), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n754), .B2(G1961), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT94), .B(G28), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(KEYINPUT30), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(new_n714), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n762), .B1(new_n764), .B2(new_n766), .C1(new_n642), .C2(new_n714), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G2084), .B2(new_n759), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n752), .A2(new_n755), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n714), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n714), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT88), .Z(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n625), .B2(new_n698), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n769), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n749), .A2(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n714), .A2(G33), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT25), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G139), .B2(new_n490), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT90), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(new_n466), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n782), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2072), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT91), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n698), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT23), .Z(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n698), .A2(G19), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT89), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n557), .B2(new_n698), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1341), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n791), .B2(new_n790), .ZN(new_n802));
  INV_X1    g377(.A(G35), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n803), .A2(KEYINPUT96), .A3(G29), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT96), .B1(new_n803), .B2(G29), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(G162), .C2(new_n714), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT29), .B(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n714), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n485), .A2(G128), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n490), .B2(G140), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(G29), .ZN(new_n817));
  INV_X1    g392(.A(G2067), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n793), .A2(new_n797), .A3(new_n802), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n748), .A2(G1996), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n781), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n736), .A2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n736), .A2(new_n823), .ZN(G150));
  NOR2_X1   g400(.A1(new_n625), .A2(new_n619), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n530), .A2(G55), .A3(G543), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n828), .B1(new_n510), .B2(new_n829), .C1(new_n830), .C2(new_n527), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n556), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n556), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n827), .B(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n836), .A2(new_n837), .A3(G860), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n831), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  AND2_X1   g416(.A1(G162), .A2(G160), .ZN(new_n842));
  NOR2_X1   g417(.A1(G162), .A2(G160), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT97), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n642), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT97), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n845), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n816), .A2(new_n508), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n816), .A2(new_n508), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n788), .B(new_n786), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n789), .A3(new_n852), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n739), .A2(new_n745), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n855), .A2(new_n746), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n721), .B(new_n630), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n490), .A2(G142), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n466), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n485), .B2(G130), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n863), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n851), .B1(new_n862), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n862), .A2(new_n851), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n850), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n869), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n861), .A3(new_n860), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n850), .A3(new_n871), .ZN(new_n877));
  XNOR2_X1  g452(.A(KEYINPUT99), .B(G37), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n874), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n874), .B2(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n556), .A2(new_n831), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n556), .A2(new_n831), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n626), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n612), .A2(new_n619), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n832), .A2(new_n889), .A3(new_n833), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  AND3_X1   g469(.A1(G299), .A2(new_n894), .A3(new_n612), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(G299), .B2(new_n612), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(G299), .B2(new_n612), .ZN(new_n899));
  AOI22_X1  g474(.A1(new_n569), .A2(new_n571), .B1(G651), .B2(new_n575), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n625), .A2(KEYINPUT102), .A3(new_n567), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n893), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n616), .A2(new_n625), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n904), .B(new_n905), .C1(new_n895), .C2(new_n896), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n892), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g483(.A1(G299), .A2(new_n612), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT101), .ZN(new_n910));
  NAND3_X1  g485(.A1(G299), .A2(new_n612), .A3(new_n894), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n910), .A2(new_n911), .B1(new_n616), .B2(new_n625), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n891), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n908), .B1(new_n907), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g490(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n703), .A2(new_n731), .ZN(new_n918));
  XNOR2_X1  g493(.A(G303), .B(G288), .ZN(new_n919));
  NAND2_X1  g494(.A1(G305), .A2(G290), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n920), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n927), .A2(new_n921), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n914), .B1(new_n915), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n930), .ZN(new_n933));
  NOR4_X1   g508(.A1(new_n933), .A2(new_n907), .A3(new_n908), .A4(new_n913), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n831), .A2(new_n621), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n885), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n899), .A2(new_n901), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n910), .A2(new_n911), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT41), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n906), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n891), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n913), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(KEYINPUT105), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n942), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n933), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n914), .A2(new_n915), .A3(new_n931), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n621), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n936), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(KEYINPUT106), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n937), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(new_n935), .A2(new_n936), .ZN(G331));
  OAI21_X1  g527(.A(G171), .B1(new_n886), .B2(new_n887), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n832), .A2(G301), .A3(new_n833), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(G168), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G168), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n897), .A2(new_n902), .A3(new_n893), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n954), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G286), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n905), .A3(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n939), .A2(new_n904), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n958), .A2(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n922), .A2(new_n923), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n878), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n961), .B2(new_n955), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n940), .A2(new_n941), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  INV_X1    g544(.A(new_n965), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G37), .B1(new_n969), .B2(new_n970), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n968), .A2(new_n958), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n975), .B2(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT43), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT44), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n966), .A2(new_n971), .A3(KEYINPUT43), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n982), .ZN(G397));
  NAND2_X1  g558(.A1(new_n816), .A2(G2067), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n811), .A2(new_n818), .A3(new_n815), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n986), .A2(new_n987), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n746), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n465), .A2(new_n501), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n504), .A2(new_n506), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n993), .A2(KEYINPUT4), .B1(new_n994), .B2(new_n479), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n494), .A2(new_n498), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n482), .A2(G2105), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n467), .A2(new_n472), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(G40), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  NOR2_X1   g579(.A1(new_n989), .A2(new_n990), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n991), .B(new_n1004), .C1(new_n1005), .C2(G1996), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1003), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(G1996), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n859), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n721), .B(new_n725), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1986), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n731), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n731), .A2(new_n1014), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1007), .B1(new_n1015), .B2(KEYINPUT107), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n1021));
  XNOR2_X1  g596(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1000), .A2(G40), .A3(new_n1001), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n998), .A2(G1384), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G114), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(KEYINPUT71), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(KEYINPUT71), .ZN(new_n1029));
  OAI21_X1  g604(.A(G2105), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(new_n496), .B1(new_n484), .B2(G126), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n499), .A2(KEYINPUT72), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n501), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n500), .B1(new_n462), .B2(new_n464), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n503), .A2(new_n1034), .B1(new_n1035), .B2(new_n499), .ZN(new_n1036));
  AOI211_X1 g611(.A(new_n1024), .B(new_n1026), .C1(new_n1031), .C2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT110), .B1(new_n508), .B2(new_n1025), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n999), .B(new_n1023), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1022), .B1(new_n1039), .B2(G2078), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1044), .A3(new_n1023), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1025), .B1(new_n995), .B2(new_n996), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n999), .A2(new_n1023), .A3(new_n773), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT53), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n508), .B2(new_n992), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1026), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1052), .A2(new_n1002), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT121), .B1(new_n1054), .B2(new_n773), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1040), .B(new_n1047), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G171), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT123), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1059), .A3(G171), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1040), .A2(G301), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1048), .A2(new_n1024), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1053), .A2(KEYINPUT110), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1052), .A2(new_n1002), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(KEYINPUT53), .A4(new_n773), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1047), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1062), .B1(new_n1063), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1068), .A2(new_n1047), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1067), .A3(new_n773), .ZN(new_n1072));
  AOI21_X1  g647(.A(G171), .B1(new_n1072), .B2(new_n1022), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT124), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1021), .B1(new_n1061), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1066), .A2(new_n1067), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  OAI211_X1 g654(.A(G40), .B(G160), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1085));
  NAND3_X1  g660(.A1(G299), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n900), .A2(KEYINPUT115), .A3(new_n1083), .A4(new_n567), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1078), .A2(new_n1082), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1078), .A2(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1045), .A2(new_n778), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1023), .A2(new_n818), .A3(new_n1042), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n625), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n1088), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT61), .B1(new_n1089), .B2(KEYINPUT118), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n625), .B(KEYINPUT119), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n612), .A2(KEYINPUT119), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1042), .A2(G160), .A3(G40), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(G1341), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1110), .A2(KEYINPUT117), .A3(new_n1112), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1115), .B(new_n1116), .C1(G1996), .C2(new_n1039), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n557), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(KEYINPUT59), .A3(new_n557), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1096), .A2(KEYINPUT61), .A3(new_n1088), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1093), .B1(new_n1109), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1073), .B(new_n1047), .C1(new_n1055), .C2(new_n1051), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1040), .ZN(new_n1126));
  OAI21_X1  g701(.A(G171), .B1(new_n1126), .B2(new_n1069), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1127), .A3(KEYINPUT54), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT125), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .A4(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n591), .A2(G1981), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT113), .B(G1981), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(KEYINPUT49), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(G8), .A3(new_n1110), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT49), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT114), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1138), .ZN(new_n1140));
  INV_X1    g715(.A(G8), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1023), .B2(new_n1042), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .A4(new_n1136), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT112), .ZN(new_n1146));
  INV_X1    g721(.A(G1976), .ZN(new_n1147));
  OR2_X1    g722(.A1(G288), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n1110), .A3(G8), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(G288), .B2(new_n1147), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1142), .A2(KEYINPUT112), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(KEYINPUT52), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1145), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(G303), .A2(G8), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT55), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G1971), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT111), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1160), .A2(new_n1161), .B1(G2090), .B2(new_n1045), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  OAI211_X1 g738(.A(G8), .B(new_n1159), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1045), .A2(G2090), .ZN(new_n1165));
  OAI21_X1  g740(.A(G8), .B1(new_n1165), .B2(new_n1160), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1158), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1156), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT51), .ZN(new_n1169));
  AND2_X1   g744(.A1(KEYINPUT120), .A2(G8), .ZN(new_n1170));
  OAI22_X1  g745(.A1(G2084), .A2(new_n1045), .B1(new_n1054), .B2(G1966), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1169), .B(new_n1170), .C1(new_n1171), .C2(G286), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(G8), .A3(G286), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g749(.A(G168), .B1(new_n1054), .B2(G1966), .C1(G2084), .C2(new_n1045), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1169), .B1(new_n1175), .B2(new_n1170), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  AND4_X1   g753(.A1(new_n1076), .A2(new_n1124), .A3(new_n1132), .A4(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1171), .A2(G8), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(G286), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1156), .A2(new_n1164), .A3(new_n1167), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(G8), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1158), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1180), .A2(new_n1183), .A3(G286), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1186), .A2(new_n1156), .A3(new_n1164), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1164), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1145), .ZN(new_n1191));
  OR2_X1    g766(.A1(G288), .A2(G1976), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1135), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1190), .A2(new_n1156), .B1(new_n1193), .B2(new_n1142), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1156), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1195));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1175), .A2(new_n1170), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT51), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1198), .A2(new_n1199), .A3(new_n1173), .A4(new_n1172), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1195), .A2(new_n1061), .A3(new_n1196), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1189), .A2(new_n1194), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1020), .B1(new_n1179), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1017), .A2(new_n1007), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT48), .Z(new_n1205));
  NAND3_X1  g780(.A1(new_n1010), .A2(new_n1012), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n991), .A2(new_n1004), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n1004), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1206), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1004), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1010), .A2(new_n722), .A3(new_n724), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n1217), .B2(new_n985), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1203), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g795(.A(G319), .B1(new_n660), .B2(new_n661), .ZN(new_n1222));
  OR2_X1    g796(.A1(G227), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g797(.A1(G229), .A2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g798(.A(new_n1224), .B1(new_n874), .B2(new_n879), .ZN(new_n1225));
  NOR2_X1   g799(.A1(new_n980), .A2(new_n981), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  OAI221_X1 g801(.A(new_n1224), .B1(new_n874), .B2(new_n879), .C1(new_n980), .C2(new_n981), .ZN(G225));
endmodule


