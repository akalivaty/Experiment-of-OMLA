//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n643, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n468), .B2(G101), .ZN(new_n469));
  AND4_X1   g044(.A1(new_n466), .A2(new_n463), .A3(G101), .A4(G2104), .ZN(new_n470));
  OAI22_X1  g045(.A1(new_n464), .A2(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n463), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n479), .B1(new_n483), .B2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n464), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n491), .B(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(KEYINPUT73), .A2(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT73), .A2(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G2105), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n462), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n500), .B(new_n501), .C1(new_n480), .C2(new_n481), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n507), .B(new_n508), .C1(new_n481), .C2(new_n480), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n508), .B1(new_n462), .B2(new_n507), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n505), .A2(new_n512), .ZN(G164));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR3_X1    g100(.A1(new_n519), .A2(new_n525), .A3(KEYINPUT74), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n519), .B2(new_n525), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n529), .A2(new_n534), .A3(G63), .A4(G651), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n521), .B2(new_n541), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n543), .A2(new_n544), .B1(G51), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n538), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  NAND3_X1  g126(.A1(new_n529), .A2(new_n534), .A3(G64), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n518), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT78), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n546), .A2(new_n547), .B1(new_n514), .B2(new_n515), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G90), .B1(new_n548), .B2(G52), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n557), .A2(G81), .B1(new_n548), .B2(G43), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n529), .A2(new_n534), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  NAND4_X1  g145(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND4_X1  g148(.A1(G319), .A2(G483), .A3(G661), .A4(new_n573), .ZN(G188));
  NAND3_X1  g149(.A1(new_n548), .A2(KEYINPUT80), .A3(G53), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n532), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n557), .A2(G91), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G166), .ZN(G303));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n518), .B1(new_n565), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G87), .ZN(new_n589));
  INV_X1    g164(.A(G49), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n521), .A2(new_n589), .B1(new_n523), .B2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n588), .A2(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(new_n548), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n557), .B2(G86), .ZN(new_n595));
  AND4_X1   g170(.A1(new_n594), .A2(new_n516), .A3(new_n520), .A4(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(G61), .B1(new_n530), .B2(new_n531), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n600), .B(G61), .C1(new_n530), .C2(new_n531), .ZN(new_n601));
  NAND2_X1  g176(.A1(G73), .A2(G543), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT82), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n598), .A2(KEYINPUT81), .B1(G73), .B2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n518), .B1(new_n606), .B2(new_n601), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n597), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G305));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  INV_X1    g187(.A(G47), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n521), .A2(new_n612), .B1(new_n523), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  INV_X1    g190(.A(G72), .ZN(new_n616));
  OAI22_X1  g191(.A1(new_n565), .A2(new_n615), .B1(new_n616), .B2(new_n545), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n518), .B1(new_n617), .B2(KEYINPUT84), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n619), .B1(new_n616), .B2(new_n545), .C1(new_n565), .C2(new_n615), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n614), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G290));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT85), .B1(new_n521), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n557), .A2(new_n625), .A3(G92), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n523), .A2(KEYINPUT86), .ZN(new_n630));
  INV_X1    g205(.A(G54), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n523), .B2(KEYINPUT86), .ZN(new_n632));
  NAND2_X1  g207(.A1(G79), .A2(G543), .ZN(new_n633));
  INV_X1    g208(.A(G66), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n532), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n630), .A2(new_n632), .B1(G651), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n624), .A2(new_n626), .A3(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G171), .B2(new_n639), .ZN(G284));
  OAI21_X1  g216(.A(new_n640), .B1(G171), .B2(new_n639), .ZN(G321));
  NAND2_X1  g217(.A1(G299), .A2(new_n639), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G168), .B2(new_n639), .ZN(G297));
  OAI21_X1  g219(.A(new_n643), .B1(G168), .B2(new_n639), .ZN(G280));
  AND3_X1   g220(.A1(new_n629), .A2(new_n636), .A3(new_n637), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT87), .B(G559), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(G860), .B2(new_n647), .ZN(G148));
  NOR2_X1   g223(.A1(new_n569), .A2(G868), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n649), .B1(G868), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT88), .ZN(G323));
  XOR2_X1   g227(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n653));
  XNOR2_X1  g228(.A(G323), .B(new_n653), .ZN(G282));
  NAND2_X1  g229(.A1(new_n462), .A2(new_n468), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2100), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n486), .A2(new_n488), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G135), .ZN(new_n662));
  OAI21_X1  g237(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n663));
  INV_X1    g238(.A(G111), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n664), .B2(G2105), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n483), .B2(G123), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(G2096), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n659), .A2(G2100), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(G2096), .ZN(new_n670));
  NAND4_X1  g245(.A1(new_n660), .A2(new_n668), .A3(new_n669), .A4(new_n670), .ZN(G156));
  INV_X1    g246(.A(KEYINPUT14), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2427), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2430), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT15), .B(G2435), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n675), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2451), .B(G2454), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT16), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1341), .B(G1348), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n677), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2443), .B(G2446), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G14), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n685), .A2(KEYINPUT91), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT91), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G401));
  XOR2_X1   g265(.A(G2084), .B(G2090), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT92), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2072), .B(G2078), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n693), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n694), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n693), .A2(new_n694), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n701), .A2(new_n692), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n692), .A2(new_n700), .A3(new_n699), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n697), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G2096), .B(G2100), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G227));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(G1971), .B(G1976), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT19), .ZN(new_n711));
  XOR2_X1   g286(.A(G1956), .B(G2474), .Z(new_n712));
  XOR2_X1   g287(.A(G1961), .B(G1966), .Z(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n712), .A2(new_n713), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n711), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n711), .A2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT20), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n720), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(G1991), .B(G1996), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n720), .B2(new_n722), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(new_n725), .B2(new_n728), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n709), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n731), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n733), .A2(new_n729), .A3(new_n708), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n732), .A2(new_n734), .ZN(G229));
  NOR2_X1   g310(.A1(G29), .A2(G35), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G162), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT29), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2090), .Z(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  INV_X1    g315(.A(G34), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G160), .B2(new_n740), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT100), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G5), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G171), .B2(new_n749), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n746), .A2(new_n747), .B1(new_n751), .B2(G1961), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(G1961), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n748), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n739), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G4), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n646), .B2(G16), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(G1348), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n463), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n661), .A2(G139), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT98), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n765), .C1(new_n759), .C2(new_n761), .ZN(new_n766));
  MUX2_X1   g341(.A(G33), .B(new_n766), .S(G29), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2072), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G168), .A2(new_n749), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n749), .B2(G21), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n758), .B(new_n768), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G32), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT102), .B1(new_n740), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G105), .B2(new_n468), .ZN(new_n778));
  INV_X1    g353(.A(G129), .ZN(new_n779));
  INV_X1    g354(.A(new_n483), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G141), .B2(new_n661), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  MUX2_X1   g358(.A(KEYINPUT102), .B(new_n774), .S(new_n783), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT27), .B(G1996), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT103), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n749), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n569), .B2(new_n749), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT96), .B(G1341), .Z(new_n789));
  OAI22_X1  g364(.A1(new_n784), .A2(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n740), .A2(G27), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G164), .B2(new_n740), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G2078), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT30), .B(G28), .ZN(new_n795));
  OR2_X1    g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  NAND2_X1  g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n795), .A2(new_n740), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n794), .B(new_n798), .C1(new_n740), .C2(new_n667), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n757), .A2(G1348), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n771), .B2(new_n769), .ZN(new_n801));
  NOR4_X1   g376(.A1(new_n790), .A2(new_n793), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n749), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  INV_X1    g379(.A(G299), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n749), .ZN(new_n806));
  INV_X1    g381(.A(G1956), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n788), .A2(new_n789), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n740), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT28), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G116), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n483), .B2(G128), .ZN(new_n816));
  INV_X1    g391(.A(G140), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n489), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n812), .B1(new_n820), .B2(new_n740), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2067), .ZN(new_n822));
  AOI211_X1 g397(.A(new_n810), .B(new_n822), .C1(new_n786), .C2(new_n784), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n755), .A2(new_n772), .A3(new_n802), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n749), .A2(G23), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n588), .A2(new_n591), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n749), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT33), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n830), .B(new_n826), .C1(new_n827), .C2(new_n749), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1976), .ZN(new_n833));
  NOR2_X1   g408(.A1(G6), .A2(G16), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n610), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT32), .B(G1981), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n835), .B(new_n836), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n749), .A2(G22), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n749), .ZN(new_n839));
  INV_X1    g414(.A(G1971), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n833), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT34), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n749), .A2(G24), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n621), .B2(new_n749), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(G1986), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n740), .A2(G25), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n661), .A2(G131), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G107), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(G2105), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n483), .B2(G119), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n847), .B1(new_n854), .B2(new_n740), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G1991), .Z(new_n856));
  XOR2_X1   g431(.A(new_n855), .B(new_n856), .Z(new_n857));
  AND2_X1   g432(.A1(new_n845), .A2(G1986), .ZN(new_n858));
  NOR4_X1   g433(.A1(new_n843), .A2(new_n846), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n842), .A2(KEYINPUT34), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n842), .A2(KEYINPUT95), .A3(KEYINPUT34), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n825), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n825), .A3(new_n864), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n824), .B1(new_n866), .B2(new_n867), .ZN(G311));
  AND3_X1   g443(.A1(new_n802), .A2(new_n772), .A3(new_n823), .ZN(new_n869));
  INV_X1    g444(.A(new_n867), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n869), .B(new_n755), .C1(new_n870), .C2(new_n865), .ZN(G150));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n872));
  XNOR2_X1  g447(.A(KEYINPUT105), .B(G860), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  INV_X1    g449(.A(G55), .ZN(new_n875));
  OAI22_X1  g450(.A1(new_n521), .A2(new_n874), .B1(new_n523), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(G80), .A2(G543), .ZN(new_n877));
  INV_X1    g452(.A(G67), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n565), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n879), .B2(G651), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n569), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n563), .A2(new_n568), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g459(.A(KEYINPUT104), .B(new_n876), .C1(new_n879), .C2(G651), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT38), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n646), .A2(G559), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n873), .B1(new_n896), .B2(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n884), .A2(new_n885), .ZN(new_n903));
  INV_X1    g478(.A(new_n873), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT107), .Z(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT37), .Z(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n872), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n901), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(new_n899), .ZN(new_n911));
  OAI211_X1 g486(.A(KEYINPUT108), .B(new_n907), .C1(new_n911), .C2(new_n897), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(G145));
  INV_X1    g488(.A(new_n781), .ZN(new_n914));
  INV_X1    g489(.A(G141), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n915), .B2(new_n489), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n916), .A2(new_n766), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n766), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n853), .B(new_n656), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n501), .B1(new_n480), .B2(new_n481), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT72), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n925), .A2(new_n503), .B1(new_n496), .B2(new_n498), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n507), .B1(new_n480), .B2(new_n481), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT4), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n509), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT109), .B1(new_n928), .B2(new_n509), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n820), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n661), .A2(G142), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT110), .Z(new_n934));
  NAND2_X1  g509(.A1(new_n483), .A2(G130), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n936), .A2(new_n463), .A3(G118), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n463), .B2(G118), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n938), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n934), .B(new_n935), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n932), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n932), .A2(new_n940), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n922), .A2(new_n923), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(G160), .B(new_n667), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(G162), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n932), .A2(new_n940), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n932), .A2(new_n940), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n916), .B(new_n766), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n921), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n943), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n945), .B1(new_n943), .B2(new_n950), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT40), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n955), .B(new_n956), .ZN(G395));
  XNOR2_X1  g532(.A(new_n887), .B(new_n650), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n646), .A2(G299), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n805), .A2(new_n638), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT112), .B1(new_n646), .B2(G299), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT41), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT41), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n961), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n958), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT42), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n526), .A2(G288), .A3(new_n527), .ZN(new_n972));
  AOI21_X1  g547(.A(G288), .B1(new_n526), .B2(new_n527), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G290), .A2(new_n610), .ZN(new_n975));
  NAND2_X1  g550(.A1(G305), .A2(new_n621), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n965), .B(new_n981), .C1(new_n958), .C2(new_n969), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n971), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n971), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(G868), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n903), .A2(new_n639), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(G295));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n986), .ZN(G331));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  NAND2_X1  g564(.A1(G286), .A2(G171), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n538), .B(new_n549), .C1(new_n556), .C2(new_n559), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n881), .A3(new_n886), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n887), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n964), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n979), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n992), .ZN(new_n997));
  INV_X1    g572(.A(new_n964), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n967), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT41), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT113), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n997), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n998), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT114), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n996), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n966), .A2(new_n994), .A3(new_n968), .A4(new_n992), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1006), .A3(new_n979), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1005), .A2(KEYINPUT43), .A3(new_n952), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n952), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n979), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT44), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1005), .A2(new_n1009), .A3(new_n952), .A4(new_n1007), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(new_n1019), .ZN(G397));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n510), .B2(new_n511), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n928), .A2(KEYINPUT109), .A3(new_n509), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n505), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n468), .A2(G101), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT68), .ZN(new_n1028));
  INV_X1    g603(.A(new_n470), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n485), .A2(G137), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n472), .A2(new_n473), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G2105), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(G40), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n818), .B(KEYINPUT97), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G2067), .ZN(new_n1036));
  INV_X1    g611(.A(G2067), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n820), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1996), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n782), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1034), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1043), .A3(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT45), .B1(new_n931), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G40), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n471), .A2(new_n474), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT116), .B1(new_n1049), .B2(G1996), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n782), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1042), .A2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(new_n853), .B(new_n856), .Z(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1034), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G290), .A2(G1986), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(new_n1057), .B2(KEYINPUT115), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1057), .A2(KEYINPUT115), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G290), .A2(G1986), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n931), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(G8), .C1(new_n1064), .C2(G288), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n827), .B2(G1976), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1063), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(G1981), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n557), .A2(G86), .B1(new_n548), .B2(G48), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n604), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n610), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(G86), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT83), .B1(new_n521), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n557), .A2(new_n594), .A3(G86), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1077), .A2(new_n1078), .B1(G48), .B2(new_n548), .ZN(new_n1079));
  AOI211_X1 g654(.A(KEYINPUT82), .B(new_n518), .C1(new_n606), .C2(new_n601), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n608), .B1(new_n603), .B2(G651), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1071), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1073), .B1(new_n1075), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT49), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1070), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1073), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1074), .B1(new_n610), .B2(new_n1071), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1082), .A2(KEYINPUT120), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1086), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1069), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n526), .A2(G8), .A3(new_n527), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1025), .B2(G1384), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n928), .A2(new_n509), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1384), .B1(new_n926), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1033), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT118), .B(G2090), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1021), .A2(G1384), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1033), .B1(new_n931), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT117), .B1(new_n1102), .B2(KEYINPUT45), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1045), .B1(new_n505), .B2(new_n512), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n1021), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n840), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1098), .A2(new_n1115), .A3(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1099), .B1(new_n931), .B2(new_n1045), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1048), .B1(new_n1110), .B2(KEYINPUT50), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n840), .A2(new_n1113), .B1(new_n1119), .B2(new_n1105), .ZN(new_n1120));
  INV_X1    g695(.A(G8), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1097), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n926), .A2(new_n1101), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1033), .B1(new_n1123), .B2(new_n1107), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1966), .B1(new_n1026), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1048), .A2(new_n747), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G286), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1094), .A2(new_n1116), .A3(new_n1122), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1097), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1128), .A2(new_n1131), .A3(G286), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1094), .A3(new_n1116), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1138), .A2(new_n1064), .A3(new_n827), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1070), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1116), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1141), .A2(new_n1142), .B1(new_n1094), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1069), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n1138), .A2(new_n1116), .A3(new_n1122), .A4(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1104), .A2(G1961), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1113), .A2(G2078), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1107), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1048), .B1(G164), .B2(new_n1151), .ZN(new_n1152));
  OR4_X1    g727(.A1(new_n1149), .A2(new_n1046), .A3(G2078), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1155));
  NAND2_X1  g730(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1030), .A2(KEYINPUT124), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1030), .A2(KEYINPUT124), .ZN(new_n1159));
  NOR4_X1   g734(.A1(new_n474), .A2(new_n1149), .A3(new_n1047), .A4(G2078), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n931), .B2(new_n1107), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1155), .A2(new_n1156), .B1(new_n1162), .B2(new_n1026), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1154), .A2(new_n1157), .B1(new_n1150), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n548), .A2(G51), .ZN(new_n1165));
  INV_X1    g740(.A(new_n544), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(G8), .B1(new_n1168), .B2(new_n537), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT122), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT51), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1128), .A2(new_n1171), .A3(new_n1169), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1169), .B2(KEYINPUT122), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n769), .B1(new_n1046), .B2(new_n1152), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1126), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT50), .B1(new_n931), .B2(new_n1045), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1110), .A2(new_n1099), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(G8), .B(new_n1174), .C1(new_n1180), .C2(G286), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1172), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1169), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT123), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1186), .B(new_n1183), .C1(new_n1172), .C2(new_n1181), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1146), .B(new_n1164), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT57), .ZN(new_n1189));
  XNOR2_X1  g764(.A(G299), .B(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n807), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1191));
  XNOR2_X1  g766(.A(KEYINPUT56), .B(G2072), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1196));
  AOI21_X1  g771(.A(G1348), .B1(new_n1196), .B2(new_n1048), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1063), .A2(G2067), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n646), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1190), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1195), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT60), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1205));
  OAI221_X1 g780(.A(KEYINPUT60), .B1(G2067), .B2(new_n1063), .C1(new_n1104), .C2(G1348), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n646), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1190), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1195), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1202), .A2(KEYINPUT61), .A3(new_n1194), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1207), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1206), .A2(new_n646), .ZN(new_n1213));
  XOR2_X1   g788(.A(KEYINPUT58), .B(G1341), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1063), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(new_n1113), .B2(G1996), .ZN(new_n1216));
  AND3_X1   g791(.A1(new_n1216), .A2(KEYINPUT59), .A3(new_n569), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT59), .B1(new_n1216), .B2(new_n569), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1213), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1203), .B1(new_n1212), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g795(.A(new_n1137), .B(new_n1144), .C1(new_n1188), .C2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1146), .A2(G171), .A3(new_n1154), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1223), .A2(new_n1186), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1182), .A2(KEYINPUT123), .A3(new_n1184), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1224), .A2(KEYINPUT62), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1227), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1222), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1062), .B1(new_n1221), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT46), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1044), .A2(new_n1050), .A3(new_n1231), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1232), .B(KEYINPUT125), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1036), .A2(new_n1038), .A3(new_n782), .ZN(new_n1234));
  AOI22_X1  g809(.A1(KEYINPUT46), .A2(new_n1051), .B1(new_n1234), .B2(new_n1034), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT47), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1233), .A2(KEYINPUT47), .A3(new_n1235), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1060), .A2(new_n1034), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1242), .B(KEYINPUT48), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n854), .A2(new_n856), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1038), .B1(new_n1053), .B2(new_n1244), .ZN(new_n1245));
  AOI22_X1  g820(.A1(new_n1055), .A2(new_n1243), .B1(new_n1245), .B2(new_n1034), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1239), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1248));
  NOR2_X1   g823(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1230), .A2(new_n1249), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g825(.A1(G227), .A2(new_n460), .ZN(new_n1252));
  AOI21_X1  g826(.A(new_n1252), .B1(new_n688), .B2(new_n687), .ZN(new_n1253));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1254));
  AOI22_X1  g828(.A1(new_n1253), .A2(new_n1254), .B1(new_n732), .B2(new_n734), .ZN(new_n1255));
  OAI21_X1  g829(.A(KEYINPUT127), .B1(G401), .B2(new_n1252), .ZN(new_n1256));
  AND2_X1   g830(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OR2_X1    g831(.A1(new_n953), .A2(new_n954), .ZN(new_n1258));
  AND3_X1   g832(.A1(new_n1257), .A2(new_n1258), .A3(new_n1017), .ZN(G308));
  NAND3_X1  g833(.A1(new_n1257), .A2(new_n1258), .A3(new_n1017), .ZN(G225));
endmodule


