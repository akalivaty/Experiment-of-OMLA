//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT22), .ZN(new_n208));
  INV_X1    g007(.A(G211gat), .ZN(new_n209));
  INV_X1    g008(.A(G218gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n207), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT29), .B1(new_n213), .B2(KEYINPUT86), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n211), .ZN(new_n215));
  INV_X1    g014(.A(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n218), .A3(new_n212), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT3), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT80), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(G155gat), .A3(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n222), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G141gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G148gat), .ZN(new_n230));
  INV_X1    g029(.A(G148gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n223), .A2(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT81), .B1(new_n231), .B2(G141gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n229), .A3(G148gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n238), .A3(new_n232), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n221), .B1(new_n227), .B2(KEYINPUT2), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n228), .A2(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n220), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n212), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n205), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT3), .B1(new_n243), .B2(new_n246), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n249), .B(new_n204), .C1(new_n241), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT87), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT31), .B(G50gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(G22gat), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G22gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n250), .A2(new_n241), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n259), .A2(new_n247), .A3(new_n205), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n249), .B1(new_n241), .B2(new_n220), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n205), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n258), .B(new_n255), .C1(new_n262), .C2(KEYINPUT87), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(KEYINPUT87), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n257), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n257), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G227gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(new_n203), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G134gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT69), .B(G134gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(new_n270), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT70), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n275), .B1(new_n277), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT71), .B1(new_n276), .B2(G120gat), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n282), .A2(new_n284), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT28), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT27), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G183gat), .ZN(new_n299));
  AND4_X1   g098(.A1(KEYINPUT28), .A2(new_n297), .A3(new_n299), .A4(new_n294), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n295), .A2(new_n300), .B1(new_n296), .B2(new_n294), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n303), .A2(KEYINPUT68), .A3(new_n306), .A4(new_n304), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n302), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n302), .B2(new_n304), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n313), .A2(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n301), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n294), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(KEYINPUT64), .A3(new_n324), .A4(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n326));
  INV_X1    g125(.A(G169gat), .ZN(new_n327));
  INV_X1    g126(.A(G176gat), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT23), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n312), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n322), .A2(new_n325), .A3(new_n326), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n303), .A2(KEYINPUT23), .A3(new_n306), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n333), .A2(KEYINPUT25), .A3(new_n330), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n321), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n331), .A2(new_n332), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n292), .B1(new_n317), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n332), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(new_n338), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n311), .A2(new_n316), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n293), .A2(new_n294), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n348), .B1(G183gat), .B2(G190gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n288), .A2(new_n291), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n273), .A2(new_n283), .A3(new_n280), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n283), .B1(new_n273), .B2(new_n280), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n269), .B1(new_n340), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT34), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT75), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n340), .A2(new_n355), .A3(new_n269), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT74), .ZN(new_n365));
  XOR2_X1   g164(.A(G71gat), .B(G99gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n362), .B(KEYINPUT32), .C1(new_n363), .C2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n369));
  NAND2_X1  g168(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n361), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n362), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT73), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n374), .A3(new_n363), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n367), .B1(new_n362), .B2(KEYINPUT32), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n340), .A2(new_n355), .ZN(new_n380));
  INV_X1    g179(.A(new_n269), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n380), .A2(new_n381), .A3(new_n369), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT76), .B1(new_n382), .B2(new_n360), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n370), .B(new_n384), .C1(new_n356), .C2(new_n359), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n267), .A2(new_n378), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n391), .B(KEYINPUT78), .Z(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n317), .B2(new_n339), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n343), .B2(new_n350), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n243), .B(new_n393), .C1(new_n394), .C2(new_n392), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(KEYINPUT79), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n397), .B(new_n392), .C1(new_n317), .C2(new_n339), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n246), .B1(new_n317), .B2(new_n339), .ZN(new_n399));
  INV_X1    g198(.A(new_n392), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n396), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n390), .B(new_n395), .C1(new_n401), .C2(new_n243), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n400), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n400), .B1(new_n343), .B2(new_n350), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n397), .ZN(new_n407));
  INV_X1    g206(.A(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n243), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n411), .A2(KEYINPUT30), .A3(new_n390), .A4(new_n395), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n395), .B1(new_n401), .B2(new_n243), .ZN(new_n413));
  INV_X1    g212(.A(new_n390), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n404), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT0), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n241), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n354), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n241), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n426), .B(KEYINPUT82), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n422), .A2(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n354), .A2(new_n431), .A3(new_n245), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n427), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n428), .B(new_n430), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT85), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n442), .A3(KEYINPUT4), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n292), .A2(new_n241), .A3(new_n433), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n432), .A2(new_n435), .A3(new_n429), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n421), .B1(new_n439), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT6), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n439), .A2(new_n448), .ZN(new_n452));
  INV_X1    g251(.A(new_n421), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n450), .B1(new_n454), .B2(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n417), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT35), .B1(new_n387), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n371), .A2(new_n458), .A3(new_n377), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n361), .A2(new_n368), .A3(new_n370), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT77), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n361), .A2(new_n370), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n379), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n449), .A2(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT88), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n448), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n453), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n439), .A2(new_n448), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT6), .B1(new_n472), .B2(new_n421), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT35), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n466), .A2(new_n475), .A3(new_n417), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n435), .B1(new_n445), .B2(new_n432), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT39), .B1(new_n425), .B2(new_n427), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT39), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(KEYINPUT40), .A3(new_n421), .A4(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n421), .B1(new_n479), .B2(new_n480), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT39), .B(new_n435), .C1(new_n445), .C2(new_n432), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n416), .A2(new_n484), .A3(new_n471), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n267), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n405), .A2(new_n393), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT37), .B1(new_n491), .B2(new_n243), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n396), .A2(new_n398), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n410), .B1(new_n493), .B2(new_n405), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT89), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n406), .B1(new_n399), .B2(new_n400), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n410), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n498), .B(new_n499), .C1(new_n410), .C2(new_n401), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT38), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  INV_X1    g301(.A(new_n395), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n409), .B2(new_n410), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n390), .B1(new_n504), .B2(new_n496), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n502), .B1(new_n501), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n414), .B1(new_n413), .B2(KEYINPUT37), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT38), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n474), .A2(new_n512), .A3(new_n402), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n490), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n267), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n456), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n386), .B2(new_n378), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n459), .A2(new_n462), .A3(new_n464), .A4(new_n517), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n478), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G57gat), .B(G64gat), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G57gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G64gat), .ZN(new_n530));
  INV_X1    g329(.A(G64gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G57gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n527), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(new_n270), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543));
  XNOR2_X1  g342(.A(G15gat), .B(G22gat), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n258), .A2(G15gat), .ZN(new_n546));
  INV_X1    g345(.A(G15gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n546), .B(new_n548), .C1(new_n549), .C2(G1gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(G8gat), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n548), .ZN(new_n553));
  INV_X1    g352(.A(G1gat), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT92), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G8gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n550), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n528), .A2(new_n536), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(KEYINPUT21), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n542), .B(new_n560), .Z(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n225), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  OR2_X1    g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(G43gat), .A2(G50gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(G43gat), .A2(G50gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT15), .B1(new_n575), .B2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n577));
  INV_X1    g376(.A(G29gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n580));
  AOI21_X1  g379(.A(G36gat), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n574), .B(new_n576), .C1(new_n581), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G36gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n580), .ZN(new_n586));
  NOR2_X1   g385(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT15), .A4(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n558), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n553), .A2(new_n554), .ZN(new_n598));
  AND4_X1   g397(.A1(new_n543), .A2(new_n598), .A3(new_n556), .A4(new_n550), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n556), .B1(new_n555), .B2(new_n550), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n591), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n584), .A2(KEYINPUT17), .A3(new_n590), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(new_n558), .B2(new_n591), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(new_n603), .A3(new_n606), .A4(new_n604), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n597), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n596), .B1(new_n610), .B2(KEYINPUT18), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n612), .B(new_n597), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT91), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G197gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT11), .B(G169gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT91), .B(new_n620), .C1(new_n611), .C2(new_n613), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G99gat), .B(G106gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(KEYINPUT8), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(G92gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT97), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(G92gat), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G85gat), .A2(G92gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT7), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT7), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(G85gat), .A3(G92gat), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g446(.A1(new_n631), .A2(new_n636), .A3(new_n642), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT97), .B(G92gat), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n641), .B1(new_n644), .B2(new_n646), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n631), .B1(new_n650), .B2(new_n636), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n603), .B(new_n604), .C1(new_n648), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n648), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n653), .A2(new_n591), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n630), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n654), .A3(new_n630), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n628), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  INV_X1    g458(.A(new_n628), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n659), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n537), .B1(new_n651), .B2(new_n648), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n650), .A2(new_n631), .A3(new_n636), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n636), .A2(new_n642), .A3(new_n647), .ZN(new_n665));
  INV_X1    g464(.A(new_n631), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n559), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT98), .B(KEYINPUT10), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n559), .A2(new_n664), .A3(new_n667), .A4(KEYINPUT10), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n663), .A2(new_n668), .ZN(new_n675));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n678), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR4_X1   g485(.A1(new_n569), .A2(new_n624), .A3(new_n662), .A4(new_n686), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n522), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n455), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n416), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G8gat), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  NAND3_X1  g494(.A1(new_n688), .A2(new_n416), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n697));
  AND3_X1   g496(.A1(new_n696), .A2(KEYINPUT100), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT100), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  OAI221_X1 g498(.A(new_n693), .B1(new_n694), .B2(new_n696), .C1(new_n698), .C2(new_n699), .ZN(G1325gat));
  AOI21_X1  g499(.A(G15gat), .B1(new_n688), .B2(new_n466), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT101), .Z(new_n702));
  AND4_X1   g501(.A1(new_n517), .A2(new_n462), .A3(new_n459), .A4(new_n464), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT102), .B1(new_n703), .B2(new_n518), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n519), .A2(new_n705), .A3(new_n520), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n547), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n702), .B1(new_n688), .B2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n688), .A2(new_n515), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT103), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT43), .B(G22gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR3_X1   g512(.A1(new_n568), .A2(new_n624), .A3(new_n686), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n522), .A2(new_n662), .A3(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n455), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n522), .B2(new_n662), .ZN(new_n719));
  INV_X1    g518(.A(new_n661), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n660), .B1(new_n659), .B2(new_n655), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n658), .B2(new_n661), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n267), .B1(new_n455), .B2(new_n417), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n495), .A2(new_n500), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT38), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n505), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT90), .ZN(new_n733));
  INV_X1    g532(.A(new_n402), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n505), .A2(new_n509), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(KEYINPUT38), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n733), .A2(new_n736), .A3(new_n474), .A4(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n489), .A2(new_n267), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n729), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n707), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n728), .B1(new_n741), .B2(new_n478), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n714), .B1(new_n719), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G29gat), .B1(new_n743), .B2(new_n455), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n717), .A2(new_n744), .ZN(G1328gat));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n417), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n585), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n416), .A2(new_n585), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT46), .B1(new_n715), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n752), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n754), .B(KEYINPUT105), .C1(new_n585), .C2(new_n747), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1329gat));
  OAI21_X1  g555(.A(G43gat), .B1(new_n743), .B2(new_n707), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n465), .A2(G43gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n715), .A2(KEYINPUT107), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT107), .B1(new_n715), .B2(new_n761), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n758), .A2(KEYINPUT47), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n757), .B(new_n765), .C1(new_n715), .C2(new_n761), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n759), .A2(new_n766), .B1(new_n767), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n715), .A2(G50gat), .A3(new_n267), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(KEYINPUT109), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n515), .B(new_n714), .C1(new_n719), .C2(new_n742), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G50gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n771), .B(new_n773), .C1(KEYINPUT109), .C2(new_n770), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n772), .A2(new_n775), .A3(G50gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n772), .B2(G50gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n777), .A3(new_n770), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n778), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI22_X1  g578(.A1(new_n740), .A2(new_n707), .B1(new_n457), .B2(new_n477), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n624), .A2(new_n686), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n780), .A2(new_n569), .A3(new_n662), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n689), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n416), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT49), .B(G64gat), .Z(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT110), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n786), .B(new_n790), .C1(new_n785), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n782), .A2(new_n793), .A3(new_n466), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n704), .A2(new_n706), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n782), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n796), .B2(new_n793), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1334gat));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n515), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g600(.A1(new_n568), .A2(new_n781), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n719), .B2(new_n742), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n455), .ZN(new_n804));
  INV_X1    g603(.A(new_n686), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n741), .A2(new_n478), .ZN(new_n806));
  INV_X1    g605(.A(new_n624), .ZN(new_n807));
  INV_X1    g606(.A(new_n662), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n568), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  INV_X1    g610(.A(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n780), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n805), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n689), .A2(new_n641), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n804), .B1(new_n817), .B2(new_n818), .ZN(G1336gat));
  INV_X1    g618(.A(new_n649), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n803), .B2(new_n417), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n417), .A2(G92gat), .A3(new_n805), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n814), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n813), .A3(KEYINPUT112), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n811), .C1(new_n780), .C2(new_n812), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n828), .A3(new_n823), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n821), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n830), .B2(new_n822), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n803), .B2(new_n707), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n465), .A2(G99gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n817), .B2(new_n833), .ZN(G1338gat));
  NOR3_X1   g633(.A1(new_n267), .A2(G106gat), .A3(new_n805), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n826), .A2(new_n828), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G106gat), .B1(new_n803), .B2(new_n267), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT53), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n814), .B2(new_n835), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n840), .B2(new_n837), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(G1339gat));
  NAND2_X1  g643(.A1(new_n689), .A2(new_n417), .ZN(new_n845));
  AOI211_X1 g644(.A(KEYINPUT54), .B(new_n676), .C1(new_n670), .C2(new_n671), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n681), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n672), .A2(new_n849), .A3(new_n673), .ZN(new_n850));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n850), .B2(new_n682), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n663), .A2(new_n668), .A3(new_n669), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n671), .A2(new_n676), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n676), .B1(new_n670), .B2(new_n671), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(KEYINPUT114), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n671), .A2(new_n676), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n849), .B1(new_n858), .B2(new_n670), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n857), .B1(new_n674), .B2(new_n859), .ZN(new_n860));
  OAI22_X1  g659(.A1(new_n848), .A2(new_n851), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n854), .B2(new_n855), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n674), .A2(new_n859), .A3(new_n857), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n847), .B1(new_n846), .B2(new_n681), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n682), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n683), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n863), .A2(new_n870), .A3(new_n622), .A4(new_n623), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n592), .A2(new_n595), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n608), .A2(new_n597), .A3(new_n609), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n618), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(new_n876));
  OR3_X1    g675(.A1(new_n611), .A2(new_n621), .A3(new_n613), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n686), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n725), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n725), .A2(new_n877), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n870), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n569), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n568), .A2(new_n624), .A3(new_n808), .A4(new_n805), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n387), .B(new_n845), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(G113gat), .B1(new_n885), .B2(new_n807), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n887), .A2(new_n515), .A3(new_n465), .A4(new_n845), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n624), .A2(new_n276), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1340gat));
  AOI21_X1  g689(.A(G120gat), .B1(new_n885), .B2(new_n686), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n805), .A2(new_n274), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n888), .B2(new_n892), .ZN(G1341gat));
  NAND3_X1  g692(.A1(new_n888), .A2(G127gat), .A3(new_n568), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n896));
  AOI21_X1  g695(.A(G127gat), .B1(new_n885), .B2(new_n568), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1342gat));
  NAND2_X1  g697(.A1(new_n888), .A2(new_n662), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n808), .A2(new_n272), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n899), .A2(G134gat), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n900), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT119), .B(new_n903), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1343gat));
  NOR2_X1   g710(.A1(new_n795), .A2(new_n845), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n515), .A2(KEYINPUT57), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n871), .A2(new_n878), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n916), .A2(new_n662), .B1(new_n881), .B2(new_n880), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n569), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n884), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n917), .B2(new_n569), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n887), .B2(new_n267), .ZN(new_n924));
  AOI211_X1 g723(.A(new_n624), .B(new_n913), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n925), .B2(new_n229), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n887), .A2(new_n267), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n912), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(G141gat), .A3(new_n624), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n925), .B2(new_n229), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n931), .A3(KEYINPUT58), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  OAI221_X1 g732(.A(new_n930), .B1(KEYINPUT121), .B2(new_n933), .C1(new_n925), .C2(new_n229), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(new_n928), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n231), .A3(new_n686), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n914), .B1(new_n883), .B2(new_n884), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n662), .B1(new_n871), .B2(new_n878), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n876), .A2(new_n662), .A3(new_n877), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n881), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n569), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n267), .B1(new_n944), .B2(new_n884), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n939), .A2(new_n940), .B1(new_n945), .B2(KEYINPUT57), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n940), .A2(new_n939), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n686), .A3(new_n912), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n938), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n913), .B1(new_n922), .B2(new_n924), .ZN(new_n951));
  AOI211_X1 g750(.A(KEYINPUT59), .B(new_n231), .C1(new_n951), .C2(new_n686), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n937), .B1(new_n950), .B2(new_n952), .ZN(G1345gat));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n225), .A3(new_n568), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n951), .A2(new_n568), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n225), .ZN(G1346gat));
  AOI21_X1  g755(.A(G162gat), .B1(new_n936), .B2(new_n662), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n726), .A2(new_n226), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n951), .B2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n887), .A2(new_n515), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n455), .A2(new_n416), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT123), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(new_n465), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n964), .A2(new_n327), .A3(new_n624), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n387), .A2(new_n961), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n887), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(G169gat), .B1(new_n968), .B2(new_n807), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n965), .A2(new_n969), .ZN(G1348gat));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n328), .A3(new_n686), .ZN(new_n971));
  OAI21_X1  g770(.A(G176gat), .B1(new_n964), .B2(new_n805), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n974), .A2(KEYINPUT60), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n968), .A2(new_n293), .A3(new_n568), .ZN(new_n976));
  OAI21_X1  g775(.A(G183gat), .B1(new_n964), .B2(new_n569), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n974), .A2(KEYINPUT60), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n978), .B(new_n979), .Z(G1350gat));
  NAND3_X1  g779(.A1(new_n968), .A2(new_n294), .A3(new_n725), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n662), .A3(new_n963), .ZN(new_n982));
  XNOR2_X1  g781(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n982), .A2(G190gat), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n982), .B2(G190gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n981), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NOR2_X1   g785(.A1(new_n795), .A2(new_n961), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n927), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n807), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n795), .A2(new_n962), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n948), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n807), .A2(G197gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1352gat));
  NAND3_X1  g792(.A1(new_n948), .A2(new_n686), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G204gat), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n805), .A2(G204gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n927), .A2(new_n987), .A3(new_n996), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT62), .Z(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n995), .A2(new_n998), .A3(KEYINPUT126), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n209), .A3(new_n568), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n568), .B(new_n990), .C1(new_n946), .C2(new_n947), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g809(.A(KEYINPUT127), .B(new_n1004), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1354gat));
  AOI21_X1  g811(.A(new_n210), .B1(new_n991), .B2(new_n662), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n988), .A2(new_n210), .A3(new_n725), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1355gat));
endmodule


