//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G113gat), .B2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G113gat), .A2(G120gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n203), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G120gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n213), .A2(new_n204), .A3(new_n206), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G127gat), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(KEYINPUT69), .A3(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT70), .B(G113gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n205), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n210), .A2(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  INV_X1    g024(.A(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G183gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT24), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n232), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  XNOR2_X1  g034(.A(G183gat), .B(G190gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(new_n225), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n240), .A2(G169gat), .A3(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT23), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(KEYINPUT64), .A3(new_n242), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  INV_X1    g047(.A(new_n245), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(new_n240), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n244), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n238), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n238), .B2(new_n251), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n230), .A2(new_n232), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n245), .A2(KEYINPUT23), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n256), .A2(new_n241), .A3(new_n243), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n226), .A2(KEYINPUT27), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT27), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G183gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n262), .A3(new_n228), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n268), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n267), .A2(new_n269), .A3(KEYINPUT67), .A4(new_n264), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT26), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n245), .A2(KEYINPUT26), .ZN(new_n275));
  INV_X1    g074(.A(new_n231), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n224), .B1(new_n259), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G227gat), .ZN(new_n281));
  INV_X1    g080(.A(G233gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n205), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT70), .B(G113gat), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n284), .B(new_n209), .C1(new_n285), .C2(new_n212), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n208), .A2(new_n203), .A3(new_n209), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n214), .B2(new_n219), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n258), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n244), .A2(new_n247), .A3(new_n250), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n233), .B2(new_n237), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n292), .B2(new_n252), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n278), .B(new_n289), .C1(new_n293), .C2(new_n253), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n280), .A2(new_n283), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT33), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n299), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n294), .ZN(new_n303));
  INV_X1    g102(.A(new_n283), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(KEYINPUT34), .B(new_n283), .C1(new_n280), .C2(new_n294), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n296), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311));
  INV_X1    g110(.A(G228gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n282), .ZN(new_n313));
  OR2_X1    g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G162gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n315), .B1(new_n328), .B2(G155gat), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n314), .A2(new_n319), .A3(new_n321), .A4(new_n316), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n323), .B(new_n324), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G211gat), .A2(G218gat), .ZN(new_n334));
  OR2_X1    g133(.A1(G211gat), .A2(G218gat), .ZN(new_n335));
  AND2_X1   g134(.A1(G197gat), .A2(G204gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G197gat), .A2(G204gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n334), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n335), .A2(new_n334), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n339), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n333), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n340), .B2(new_n344), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n313), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n324), .B1(new_n349), .B2(KEYINPUT79), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n353), .B(KEYINPUT29), .C1(new_n340), .C2(new_n344), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n313), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n333), .B2(new_n346), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT80), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n351), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G78gat), .B(G106gat), .Z(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n311), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G22gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n351), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n355), .A2(new_n360), .A3(new_n357), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n360), .B1(new_n355), .B2(new_n357), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT81), .B1(new_n373), .B2(new_n366), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n373), .A2(new_n366), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n377), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n374), .A2(new_n375), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT81), .B(G22gat), .C1(new_n373), .C2(new_n366), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n294), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n238), .A2(new_n251), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT66), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n238), .A2(new_n251), .A3(new_n252), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n290), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n289), .B1(new_n387), .B2(new_n278), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT34), .B1(new_n389), .B2(new_n283), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n303), .A2(new_n302), .A3(new_n304), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT33), .B1(new_n389), .B2(new_n283), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n390), .B(new_n391), .C1(new_n392), .C2(new_n299), .ZN(new_n393));
  INV_X1    g192(.A(new_n296), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n307), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n310), .A2(new_n378), .A3(new_n382), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT74), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n289), .B2(new_n348), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT72), .B(G162gat), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT2), .B1(new_n400), .B2(new_n320), .ZN(new_n401));
  INV_X1    g200(.A(new_n330), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n401), .A2(new_n402), .B1(new_n317), .B2(new_n322), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n224), .A2(KEYINPUT74), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n289), .A2(new_n348), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT73), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n289), .A3(new_n331), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n405), .A2(new_n407), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n404), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n224), .B2(new_n403), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n289), .A2(KEYINPUT75), .A3(new_n348), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT5), .B(new_n413), .C1(new_n418), .C2(new_n410), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n399), .B1(new_n289), .B2(new_n348), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n414), .B2(KEYINPUT4), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n412), .A2(new_n423), .A3(new_n410), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(KEYINPUT76), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT76), .B1(new_n422), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n419), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT0), .ZN(new_n430));
  XNOR2_X1  g229(.A(G57gat), .B(G85gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n289), .A2(new_n348), .A3(new_n397), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT74), .B1(new_n224), .B2(new_n403), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT4), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n439), .A3(new_n420), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n425), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n432), .A3(new_n419), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n436), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n432), .B1(new_n443), .B2(new_n419), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n435), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n449), .B(new_n278), .C1(new_n293), .C2(new_n253), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n332), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n387), .B2(new_n278), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n346), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n254), .A2(new_n258), .ZN(new_n456));
  INV_X1    g255(.A(new_n277), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n270), .B2(new_n271), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n456), .A2(new_n386), .B1(new_n458), .B2(new_n273), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n450), .B(new_n345), .C1(new_n459), .C2(new_n453), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G64gat), .B(G92gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OR3_X1    g264(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n460), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n452), .B1(new_n259), .B2(new_n279), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n345), .B1(new_n468), .B2(new_n450), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n460), .A3(new_n464), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(KEYINPUT30), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n448), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT85), .B1(new_n396), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n393), .A2(new_n394), .A3(new_n307), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n394), .B1(new_n393), .B2(new_n307), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n380), .A2(new_n381), .A3(new_n379), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n377), .B1(new_n369), .B2(new_n376), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n445), .A2(new_n447), .B1(new_n466), .B2(new_n472), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n478), .A2(new_n479), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n475), .A2(KEYINPUT35), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT71), .B1(new_n476), .B2(new_n477), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n439), .A2(new_n412), .A3(new_n420), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(new_n409), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n432), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n410), .B1(new_n422), .B2(new_n412), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n416), .A2(new_n417), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n398), .A3(new_n404), .A4(new_n410), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n496), .B2(KEYINPUT39), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n494), .A3(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n446), .B1(new_n500), .B2(KEYINPUT40), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT40), .ZN(new_n502));
  INV_X1    g301(.A(new_n499), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n503), .A2(new_n493), .A3(new_n497), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n504), .B2(new_n492), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n501), .A2(new_n466), .A3(new_n472), .A4(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n464), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n461), .B2(new_n465), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n455), .B2(new_n460), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT38), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n445), .A3(new_n447), .A4(new_n471), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n455), .A2(KEYINPUT83), .A3(new_n460), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT83), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n346), .C1(new_n451), .C2(new_n454), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT37), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT84), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n508), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT38), .B1(new_n470), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n455), .A2(KEYINPUT83), .A3(new_n460), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT84), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT37), .A4(new_n515), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n517), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n482), .B(new_n506), .C1(new_n512), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n382), .A2(new_n378), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n474), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n476), .C2(new_n477), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n488), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  OAI211_X1 g328(.A(KEYINPUT85), .B(new_n529), .C1(new_n396), .C2(new_n474), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n485), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n485), .A2(new_n528), .A3(KEYINPUT86), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(G1gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(new_n540), .C1(G1gat), .C2(new_n537), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G50gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G43gat), .ZN(new_n545));
  INV_X1    g344(.A(G43gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G50gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n548), .A2(KEYINPUT87), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT15), .B1(new_n548), .B2(KEYINPUT87), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n552), .B2(KEYINPUT88), .ZN(new_n555));
  INV_X1    g354(.A(G29gat), .ZN(new_n556));
  INV_X1    g355(.A(G36gat), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n553), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n546), .B2(G50gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n547), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n545), .A2(new_n561), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n552), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n566), .A2(new_n554), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n565), .B(new_n567), .C1(new_n549), .C2(new_n550), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n559), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT17), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n571), .B1(new_n559), .B2(new_n568), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n543), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n541), .B(G8gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n569), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n575), .B(new_n569), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(new_n574), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G197gat), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT11), .B(G169gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n573), .A2(KEYINPUT18), .A3(new_n574), .A4(new_n576), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n582), .B2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n536), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT92), .A3(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  AND2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n597), .A2(KEYINPUT9), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n543), .B1(new_n596), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n608), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n596), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G127gat), .ZN(new_n616));
  XOR2_X1   g415(.A(G183gat), .B(G211gat), .Z(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(new_n618), .A3(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(G85gat), .A3(G92gat), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT7), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT7), .B1(new_n625), .B2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G99gat), .ZN(new_n635));
  INV_X1    g434(.A(G106gat), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT8), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n634), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT97), .B1(new_n634), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n630), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G99gat), .B(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n630), .B(new_n641), .C1(new_n638), .C2(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n570), .B2(new_n572), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n569), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n649));
  NAND2_X1  g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n646), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n649), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n653), .B(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n623), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n660), .A3(new_n605), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT7), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n626), .B1(G85gat), .B2(G92gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT7), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n634), .A2(KEYINPUT97), .A3(new_n637), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n670));
  INV_X1    g469(.A(new_n633), .ZN(new_n671));
  NOR2_X1   g470(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n671), .A2(new_n672), .A3(G92gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n637), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n668), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n605), .B1(new_n676), .B2(new_n641), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n641), .B(KEYINPUT98), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n640), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n605), .A2(new_n645), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT99), .B1(new_n680), .B2(new_n660), .ZN(new_n681));
  INV_X1    g480(.A(new_n644), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n675), .A2(new_n669), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n641), .B1(new_n683), .B2(new_n630), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n605), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n605), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n679), .A2(new_n686), .A3(new_n644), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n685), .A2(KEYINPUT99), .A3(new_n660), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n662), .B1(new_n681), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G230gat), .A2(G233gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n680), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n685), .A2(new_n660), .A3(new_n687), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n661), .B1(new_n702), .B2(new_n688), .ZN(new_n703));
  INV_X1    g502(.A(new_n691), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n693), .B(new_n697), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n659), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n659), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n202), .A2(new_n535), .A3(new_n595), .A4(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n595), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n533), .B2(new_n534), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n202), .B1(new_n715), .B2(new_n712), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n448), .B(KEYINPUT102), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(G1gat), .Z(G1324gat));
  INV_X1    g520(.A(new_n473), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n713), .B2(new_n716), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT103), .B(new_n722), .C1(new_n713), .C2(new_n716), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(G8gat), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT16), .B(G8gat), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n725), .B2(new_n726), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n727), .B(new_n730), .C1(new_n731), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g531(.A1(new_n488), .A2(new_n527), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G15gat), .B1(new_n717), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n478), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(G15gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n717), .B2(new_n737), .ZN(G1326gat));
  NOR2_X1   g537(.A1(new_n717), .A2(new_n482), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT43), .B(G22gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(new_n658), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n623), .A2(new_n706), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n715), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n556), .A3(new_n718), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n533), .B2(new_n534), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n531), .B2(new_n742), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n593), .A2(new_n589), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT104), .B1(new_n754), .B2(new_n719), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G29gat), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n754), .A2(KEYINPUT104), .A3(new_n719), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n746), .B1(new_n756), .B2(new_n757), .ZN(G1328gat));
  NAND3_X1  g557(.A1(new_n744), .A2(new_n557), .A3(new_n722), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n754), .B2(new_n473), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(G1329gat));
  XOR2_X1   g562(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n764));
  OAI21_X1  g563(.A(G43gat), .B1(new_n754), .B2(new_n734), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(KEYINPUT106), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n748), .A2(new_n734), .A3(new_n749), .A4(new_n752), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT106), .B1(new_n767), .B2(new_n546), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n546), .A3(new_n478), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n765), .A2(KEYINPUT47), .A3(new_n769), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1330gat));
  NOR3_X1   g572(.A1(new_n754), .A2(new_n544), .A3(new_n482), .ZN(new_n774));
  AOI21_X1  g573(.A(G50gat), .B1(new_n744), .B2(new_n525), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n774), .A2(KEYINPUT48), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(KEYINPUT48), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1331gat));
  INV_X1    g577(.A(new_n751), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n659), .A2(new_n779), .A3(new_n706), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n531), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n718), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g583(.A(new_n473), .B(KEYINPUT107), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n781), .B2(new_n734), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n736), .A2(G71gat), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n525), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g596(.A1(new_n748), .A2(new_n749), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n623), .A2(new_n751), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n706), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n631), .A2(new_n633), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n802), .A3(new_n718), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n531), .A2(new_n742), .A3(new_n799), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n707), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n802), .B1(new_n809), .B2(new_n718), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT108), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n812));
  INV_X1    g611(.A(new_n809), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n719), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n803), .B(new_n812), .C1(new_n814), .C2(new_n802), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n632), .A3(new_n785), .ZN(new_n817));
  NAND2_X1  g616(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n798), .A2(new_n786), .A3(new_n800), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n801), .A2(new_n722), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n809), .A2(new_n632), .A3(new_n785), .ZN(new_n824));
  AOI22_X1  g623(.A1(G92gat), .A2(new_n823), .B1(new_n824), .B2(KEYINPUT109), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n825), .B2(new_n820), .ZN(G1337gat));
  NOR3_X1   g625(.A1(new_n798), .A2(new_n734), .A3(new_n800), .ZN(new_n827));
  XOR2_X1   g626(.A(KEYINPUT110), .B(G99gat), .Z(new_n828));
  AND2_X1   g627(.A1(new_n807), .A2(new_n808), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n478), .A2(new_n706), .A3(new_n828), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT111), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n831), .ZN(G1338gat));
  NOR3_X1   g631(.A1(new_n798), .A2(new_n482), .A3(new_n800), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n525), .A2(new_n636), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n833), .A2(new_n636), .B1(new_n813), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  OAI221_X1 g636(.A(new_n837), .B1(new_n813), .B2(new_n834), .C1(new_n833), .C2(new_n636), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1339gat));
  INV_X1    g638(.A(new_n623), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n661), .A2(new_n691), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(new_n681), .B2(new_n689), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n702), .A2(new_n688), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n704), .B1(new_n844), .B2(new_n662), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT55), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n690), .A2(new_n847), .A3(new_n691), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n698), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n705), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n697), .B1(new_n845), .B2(new_n847), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n842), .B(KEYINPUT54), .C1(new_n703), .C2(new_n704), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT112), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n705), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n847), .B1(new_n844), .B2(new_n841), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n692), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n851), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n852), .A2(new_n698), .A3(new_n848), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n856), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n854), .A2(new_n863), .A3(new_n751), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n579), .A2(new_n581), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n574), .B1(new_n573), .B2(new_n576), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n586), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n706), .A2(new_n589), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n742), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n589), .A2(new_n867), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n658), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n854), .A2(new_n863), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n840), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n659), .A2(new_n779), .A3(new_n707), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT113), .B1(new_n875), .B2(new_n482), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n877));
  AOI211_X1 g676(.A(new_n877), .B(new_n525), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n719), .A2(new_n736), .A3(new_n785), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n714), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n719), .B1(new_n873), .B2(new_n874), .ZN(new_n883));
  INV_X1    g682(.A(new_n396), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n786), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n285), .A3(new_n751), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n882), .A2(new_n887), .ZN(G1340gat));
  AOI21_X1  g687(.A(G120gat), .B1(new_n886), .B2(new_n706), .ZN(new_n889));
  INV_X1    g688(.A(new_n881), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n707), .A2(new_n212), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n881), .B2(new_n840), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n886), .A2(new_n217), .A3(new_n623), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1342gat));
  NOR2_X1   g694(.A1(new_n722), .A2(new_n658), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n885), .A2(new_n215), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT56), .Z(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n881), .B2(new_n658), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n733), .A2(new_n482), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n901), .ZN(new_n902));
  NOR4_X1   g701(.A1(new_n902), .A2(G141gat), .A3(new_n714), .A4(new_n785), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n733), .A2(new_n719), .A3(new_n785), .ZN(new_n907));
  XOR2_X1   g706(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(new_n875), .B2(new_n525), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n525), .A2(KEYINPUT57), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n861), .A2(KEYINPUT115), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n853), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n911), .A2(new_n595), .A3(new_n913), .A4(new_n859), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n742), .B1(new_n914), .B2(new_n868), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n840), .B1(new_n915), .B2(new_n872), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n916), .B2(new_n874), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n907), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n906), .B(G141gat), .C1(new_n918), .C2(new_n714), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n905), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n918), .A2(new_n779), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n921), .A2(G141gat), .B1(new_n904), .B2(new_n903), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n906), .ZN(G1344gat));
  AND2_X1   g722(.A1(new_n883), .A2(new_n901), .ZN(new_n924));
  INV_X1    g723(.A(G148gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n706), .A4(new_n786), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT117), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n525), .A2(new_n908), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n873), .B2(new_n874), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR4_X1   g731(.A1(new_n850), .A2(new_n658), .A3(new_n853), .A4(new_n870), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n840), .B1(new_n915), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n709), .A2(new_n714), .A3(new_n711), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n482), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n929), .A2(new_n930), .B1(new_n936), .B2(KEYINPUT57), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n907), .A2(new_n706), .ZN(new_n939));
  OAI21_X1  g738(.A(G148gat), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT59), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n918), .B2(new_n707), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT118), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n943), .A2(KEYINPUT118), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n927), .B1(new_n945), .B2(new_n946), .ZN(G1345gat));
  OAI21_X1  g746(.A(G155gat), .B1(new_n918), .B2(new_n840), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n924), .A2(new_n320), .A3(new_n623), .A4(new_n786), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(G1346gat));
  OAI21_X1  g749(.A(new_n328), .B1(new_n918), .B2(new_n658), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n924), .A2(new_n400), .A3(new_n896), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1347gat));
  NOR3_X1   g752(.A1(new_n718), .A2(new_n473), .A3(new_n736), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n879), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(G169gat), .B1(new_n955), .B2(new_n714), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n718), .B1(new_n873), .B2(new_n874), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(new_n884), .A3(new_n785), .ZN(new_n960));
  INV_X1    g759(.A(G169gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(new_n961), .A3(new_n751), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT120), .Z(new_n963));
  OAI211_X1 g762(.A(KEYINPUT121), .B(G169gat), .C1(new_n955), .C2(new_n714), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n958), .A2(new_n963), .A3(new_n964), .ZN(G1348gat));
  OAI21_X1  g764(.A(G176gat), .B1(new_n955), .B2(new_n707), .ZN(new_n966));
  INV_X1    g765(.A(G176gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n960), .A2(new_n967), .A3(new_n706), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(G1349gat));
  NAND4_X1  g768(.A1(new_n960), .A2(new_n260), .A3(new_n262), .A4(new_n623), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n623), .B(new_n954), .C1(new_n876), .C2(new_n878), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(new_n226), .ZN(new_n973));
  AND2_X1   g772(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n228), .A3(new_n742), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n742), .B(new_n954), .C1(new_n876), .C2(new_n878), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n977), .A2(new_n978), .A3(G190gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(KEYINPUT123), .B(new_n976), .C1(new_n979), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1351gat));
  OAI21_X1  g784(.A(KEYINPUT124), .B1(new_n932), .B2(new_n937), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n929), .A2(new_n930), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n936), .A2(KEYINPUT57), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT124), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n931), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n734), .A2(new_n722), .A3(new_n719), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n986), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n993), .A2(new_n994), .A3(new_n714), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n733), .A2(new_n482), .A3(new_n786), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n959), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n751), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n995), .A2(new_n999), .ZN(G1352gat));
  OAI21_X1  g799(.A(G204gat), .B1(new_n993), .B2(new_n707), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n997), .A2(G204gat), .A3(new_n707), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1353gat));
  OR3_X1    g803(.A1(new_n997), .A2(G211gat), .A3(new_n840), .ZN(new_n1005));
  OAI211_X1 g804(.A(new_n623), .B(new_n992), .C1(new_n932), .C2(new_n937), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  AOI21_X1  g808(.A(G218gat), .B1(new_n998), .B2(new_n742), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT126), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n993), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n742), .A2(G218gat), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1013), .B1(new_n993), .B2(new_n1011), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1010), .B1(new_n1012), .B2(new_n1014), .ZN(G1355gat));
endmodule


