//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n953, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT71), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G15gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT1), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n212), .A2(new_n213), .A3(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(new_n215), .B2(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n213), .A2(G134gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n211), .B1(new_n218), .B2(KEYINPUT69), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT70), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n208), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(new_n210), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n215), .A2(G127gat), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n217), .A2(new_n226), .A3(KEYINPUT1), .ZN(new_n227));
  AOI22_X1  g026(.A1(new_n219), .A2(new_n221), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n237), .B2(KEYINPUT24), .ZN(new_n238));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT23), .ZN(new_n240));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT25), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n239), .B2(KEYINPUT23), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(G169gat), .A3(G176gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n247), .A2(new_n243), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G183gat), .B(G190gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n231), .B1(new_n252), .B2(new_n230), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n229), .B1(new_n245), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n246), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n248), .A2(new_n243), .A3(new_n250), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n247), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n259), .A3(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n239), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n262), .A2(KEYINPUT26), .ZN(new_n263));
  INV_X1    g062(.A(new_n241), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n262), .B2(KEYINPUT26), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n263), .A2(new_n265), .B1(G183gat), .B2(G190gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n233), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(G190gat), .B1(new_n233), .B2(KEYINPUT27), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n273), .B2(KEYINPUT67), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n268), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n276), .B(KEYINPUT28), .C1(KEYINPUT27), .C2(new_n233), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n228), .B1(new_n261), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n276), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n271), .A2(KEYINPUT27), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n285));
  OAI21_X1  g084(.A(G183gat), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT28), .B1(new_n288), .B2(new_n274), .ZN(new_n289));
  INV_X1    g088(.A(new_n279), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n266), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n218), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g091(.A(new_n211), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n221), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n227), .A2(new_n225), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n291), .A2(new_n255), .A3(new_n260), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n206), .B1(new_n299), .B2(KEYINPUT33), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n282), .B1(new_n281), .B2(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT34), .B(new_n282), .C1(new_n281), .C2(new_n297), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n206), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT33), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n298), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n301), .A2(new_n302), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(new_n304), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n306), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n308), .B1(new_n306), .B2(new_n313), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT36), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n306), .A2(new_n313), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n306), .A2(new_n308), .A3(new_n313), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT36), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT72), .B1(new_n261), .B2(new_n280), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n291), .A2(new_n327), .A3(new_n255), .A4(new_n260), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n245), .A2(new_n254), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT29), .B1(new_n291), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT73), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n280), .A2(new_n330), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n334), .B(new_n325), .C1(new_n335), .C2(KEYINPUT29), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338));
  INV_X1    g137(.A(G211gat), .ZN(new_n339));
  INV_X1    g138(.A(G218gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n333), .A3(new_n336), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n324), .A2(new_n347), .A3(new_n328), .A4(new_n325), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n335), .A2(new_n326), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT74), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n346), .A2(new_n350), .A3(new_n357), .A4(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n355), .A2(KEYINPUT75), .A3(new_n356), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  INV_X1    g164(.A(G141gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n366), .A2(G148gat), .ZN(new_n367));
  INV_X1    g166(.A(G148gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G141gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n366), .B2(G148gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(G148gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n372), .A2(new_n365), .ZN(new_n379));
  NAND2_X1  g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n370), .A2(new_n373), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n294), .A2(new_n295), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT4), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n228), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  XNOR2_X1  g189(.A(G141gat), .B(G148gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n373), .B1(new_n391), .B2(KEYINPUT2), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n389), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n388), .B1(new_n395), .B2(new_n296), .ZN(new_n396));
  NOR4_X1   g195(.A1(new_n228), .A2(new_n393), .A3(new_n394), .A4(KEYINPUT77), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n364), .B(new_n387), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n296), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n383), .ZN(new_n402));
  INV_X1    g201(.A(new_n364), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n382), .A2(new_n390), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT77), .B1(new_n408), .B2(new_n228), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n395), .A2(new_n388), .A3(new_n296), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n384), .A2(new_n386), .A3(KEYINPUT80), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n386), .A2(KEYINPUT80), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n403), .A2(KEYINPUT5), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT79), .ZN(new_n418));
  XOR2_X1   g217(.A(G57gat), .B(G85gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT81), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n424), .B(new_n425), .C1(new_n423), .C2(new_n416), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n415), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n416), .A2(new_n423), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n427), .B2(new_n422), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT81), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n426), .A2(new_n428), .A3(new_n431), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n346), .A2(new_n350), .ZN(new_n437));
  INV_X1    g236(.A(new_n353), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n356), .B2(new_n354), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n363), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n344), .A2(KEYINPUT29), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n443), .A2(KEYINPUT83), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n390), .B1(new_n443), .B2(KEYINPUT83), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n400), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n345), .B1(new_n406), .B2(new_n347), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n447), .A2(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(KEYINPUT84), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G228gat), .ZN(new_n451));
  INV_X1    g250(.A(G233gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(new_n400), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n407), .A3(new_n453), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(new_n447), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G50gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G22gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(KEYINPUT85), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n466), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n455), .A2(new_n458), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n323), .B1(new_n442), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n423), .B1(new_n427), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n416), .A2(KEYINPUT87), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n434), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n431), .A2(new_n428), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n355), .A2(new_n358), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n438), .A2(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n437), .B2(new_n438), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n329), .A2(new_n333), .A3(new_n336), .A4(new_n344), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n348), .A2(new_n345), .A3(new_n349), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT37), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT38), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n437), .A2(KEYINPUT37), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT38), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n478), .A2(new_n479), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n471), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n440), .B1(new_n361), .B2(new_n362), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n403), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(new_n423), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n403), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(KEYINPUT39), .C1(new_n403), .C2(new_n402), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT40), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT88), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT88), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n496), .A2(new_n498), .A3(new_n502), .A4(KEYINPUT40), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT86), .B(KEYINPUT40), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n499), .A2(new_n505), .B1(new_n475), .B2(new_n474), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n490), .B(new_n491), .C1(new_n492), .C2(new_n507), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n314), .A2(new_n315), .A3(new_n471), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n363), .A2(new_n509), .A3(new_n436), .A4(new_n441), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n492), .A3(new_n509), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n472), .A2(new_n508), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT96), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT13), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n463), .A2(G15gat), .ZN(new_n518));
  INV_X1    g317(.A(G15gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G22gat), .ZN(new_n520));
  INV_X1    g319(.A(G1gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT16), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G8gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n524), .C1(G1gat), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT94), .ZN(new_n527));
  AOI21_X1  g326(.A(G1gat), .B1(new_n518), .B2(new_n520), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n524), .A4(new_n523), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n524), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n523), .B(KEYINPUT92), .C1(G1gat), .C2(new_n525), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT93), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT93), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n205), .A2(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(G50gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G43gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT15), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(KEYINPUT90), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G50gat), .ZN(new_n547));
  AOI21_X1  g346(.A(G43gat), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n205), .B2(G50gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n540), .A2(KEYINPUT89), .A3(G43gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n544), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT14), .B(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G29gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n543), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n542), .B1(new_n556), .B2(new_n558), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n538), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n562), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n517), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n553), .A2(new_n559), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n542), .ZN(new_n567));
  INV_X1    g366(.A(new_n561), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT91), .A2(KEYINPUT17), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n570), .B(new_n571), .C1(new_n560), .C2(new_n561), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n538), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n532), .B(KEYINPUT95), .C1(new_n536), .C2(new_n537), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n516), .A3(new_n564), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n565), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G197gat), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT11), .B(G169gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n516), .A4(new_n564), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n582), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n514), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(G230gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n452), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT98), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G99gat), .A3(G106gat), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT8), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(KEYINPUT97), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n599), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT99), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT8), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n598), .A3(new_n608), .A4(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  INV_X1    g415(.A(G71gat), .ZN(new_n617));
  INV_X1    g416(.A(G78gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G71gat), .B(G78gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(new_n621), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(KEYINPUT99), .B(new_n599), .C1(new_n604), .C2(new_n609), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n610), .A2(new_n623), .A3(new_n624), .A4(new_n613), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT101), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n627), .A2(new_n632), .A3(new_n628), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n626), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n625), .A2(new_n628), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n597), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(new_n629), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(new_n597), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n595), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n631), .A2(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n641), .B(new_n595), .C1(new_n643), .C2(new_n597), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n625), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(G231gat), .A3(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n625), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G127gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n213), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n625), .A2(new_n647), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n538), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n662));
  INV_X1    g461(.A(G155gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n664), .B(new_n665), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n659), .A2(new_n660), .A3(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(G232gat), .A2(G233gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(KEYINPUT41), .ZN(new_n672));
  XNOR2_X1  g471(.A(G134gat), .B(G162gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n575), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(G190gat), .B(G218gat), .Z(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n635), .A2(new_n562), .B1(KEYINPUT41), .B2(new_n671), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n680), .B1(new_n678), .B2(new_n681), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n675), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n684), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n674), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n646), .A2(new_n670), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n436), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n436), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n592), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g496(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n698));
  INV_X1    g497(.A(new_n492), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n592), .A2(new_n699), .A3(new_n690), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(G8gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(KEYINPUT42), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n703), .B(new_n704), .C1(new_n700), .C2(new_n705), .ZN(G1325gat));
  NOR3_X1   g505(.A1(new_n514), .A2(new_n591), .A3(new_n689), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n314), .A2(new_n315), .ZN(new_n708));
  AOI21_X1  g507(.A(G15gat), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n323), .A2(G15gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT105), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n707), .B2(new_n711), .ZN(G1326gat));
  NAND2_X1  g511(.A1(new_n707), .A2(new_n471), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT43), .B(G22gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  NAND2_X1  g514(.A1(new_n442), .A2(new_n471), .ZN(new_n716));
  INV_X1    g515(.A(new_n323), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n508), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n511), .A2(new_n513), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n688), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n590), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n582), .A2(new_n587), .A3(new_n588), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n646), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n670), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n557), .A3(new_n695), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n514), .B2(new_n688), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n718), .A2(new_n719), .ZN(new_n732));
  INV_X1    g531(.A(new_n688), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(KEYINPUT44), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n725), .A2(new_n723), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT106), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n731), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n731), .A2(new_n734), .A3(KEYINPUT107), .A4(new_n736), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n739), .A2(new_n695), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n729), .B1(new_n557), .B2(new_n741), .ZN(G1328gat));
  NAND3_X1  g541(.A1(new_n739), .A2(new_n699), .A3(new_n740), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n739), .A2(new_n745), .A3(new_n699), .A4(new_n740), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(G36gat), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n726), .A2(G36gat), .A3(new_n492), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(new_n708), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n726), .A2(G43gat), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G43gat), .B1(new_n737), .B2(new_n717), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT47), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n323), .A3(new_n740), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(G43gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n757), .B2(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g557(.A1(new_n545), .A2(new_n547), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n726), .A2(new_n491), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n737), .B2(new_n491), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT48), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n739), .A2(new_n471), .A3(new_n740), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(new_n760), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(G1331gat));
  INV_X1    g567(.A(new_n670), .ZN(new_n769));
  NOR4_X1   g568(.A1(new_n723), .A2(new_n769), .A3(new_n733), .A4(new_n646), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n732), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n694), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g572(.A1(new_n771), .A2(new_n492), .ZN(new_n774));
  NOR2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  AND2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n774), .B2(new_n775), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n771), .B2(new_n717), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n708), .A2(new_n617), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g581(.A1(new_n771), .A2(new_n491), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n618), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n723), .A2(new_n670), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n646), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n731), .A2(new_n734), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788), .B2(new_n694), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NOR4_X1   g589(.A1(new_n514), .A2(new_n790), .A3(new_n688), .A4(new_n786), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n720), .B2(new_n785), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n694), .A2(G85gat), .A3(new_n646), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(G1336gat));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n731), .A2(new_n734), .A3(new_n699), .A4(new_n787), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n492), .A2(G92gat), .A3(new_n646), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n791), .B2(new_n792), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n800), .B(KEYINPUT110), .Z(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n791), .B2(new_n792), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n799), .B1(new_n798), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n796), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n798), .A2(new_n801), .A3(new_n799), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n720), .A2(new_n785), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n790), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n785), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n811), .A2(new_n803), .B1(new_n797), .B2(G92gat), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n807), .B(KEYINPUT111), .C1(new_n812), .C2(new_n799), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n813), .ZN(G1337gat));
  NOR2_X1   g613(.A1(new_n788), .A2(new_n717), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT112), .B(G99gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n708), .A2(new_n724), .A3(new_n816), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n815), .A2(new_n816), .B1(new_n793), .B2(new_n817), .ZN(G1338gat));
  OAI21_X1  g617(.A(G106gat), .B1(new_n788), .B2(new_n491), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n491), .A2(G106gat), .A3(new_n646), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT113), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n793), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g622(.A(new_n597), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n635), .B2(new_n636), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n634), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT55), .B1(new_n827), .B2(new_n638), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n634), .A2(new_n637), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n824), .ZN(new_n831));
  INV_X1    g630(.A(new_n595), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n644), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT115), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n826), .B(KEYINPUT54), .C1(new_n643), .C2(new_n597), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n832), .A4(new_n831), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n838), .A3(new_n644), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n833), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n835), .A2(new_n723), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n516), .B1(new_n579), .B2(new_n564), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n563), .A2(new_n564), .A3(new_n517), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n586), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n722), .B(new_n846), .C1(new_n642), .C2(new_n645), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n733), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n722), .A2(new_n685), .A3(new_n687), .A4(new_n846), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n835), .A2(new_n839), .A3(new_n842), .A4(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n769), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n769), .A2(new_n733), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n853), .A2(new_n646), .A3(KEYINPUT114), .A4(new_n591), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n689), .B2(new_n723), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n471), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n694), .A2(new_n699), .A3(new_n751), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n723), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n591), .A2(new_n209), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  AOI21_X1  g667(.A(G120gat), .B1(new_n862), .B2(new_n724), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n646), .A2(new_n207), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n866), .B2(new_n870), .ZN(G1341gat));
  NAND3_X1  g670(.A1(new_n862), .A2(new_n213), .A3(new_n670), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n769), .B1(new_n864), .B2(new_n865), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n213), .ZN(G1342gat));
  NOR3_X1   g673(.A1(new_n699), .A2(G134gat), .A3(new_n688), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n708), .A3(new_n695), .A4(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT56), .Z(new_n877));
  AOI21_X1  g676(.A(new_n688), .B1(new_n864), .B2(new_n865), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n215), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n877), .B(KEYINPUT117), .C1(new_n878), .C2(new_n215), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1343gat));
  AOI21_X1  g682(.A(new_n491), .B1(new_n852), .B2(new_n858), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n694), .A2(new_n699), .A3(new_n323), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n591), .A2(G141gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n491), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n837), .B(new_n644), .C1(new_n589), .C2(new_n590), .ZN(new_n891));
  XOR2_X1   g690(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n892));
  AOI21_X1  g691(.A(new_n595), .B1(new_n638), .B2(new_n830), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n836), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n847), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n688), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n670), .B1(new_n896), .B2(new_n850), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n890), .B1(new_n897), .B2(new_n857), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT119), .B(new_n890), .C1(new_n897), .C2(new_n857), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n852), .A2(new_n858), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT57), .B1(new_n903), .B2(new_n471), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n885), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT120), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n907), .B(new_n885), .C1(new_n902), .C2(new_n904), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n723), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n888), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n887), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n723), .B(new_n885), .C1(new_n902), .C2(new_n904), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(G141gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  AOI211_X1 g715(.A(new_n916), .B(new_n912), .C1(new_n913), .C2(G141gat), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n910), .A2(new_n911), .B1(new_n915), .B2(new_n917), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n471), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n830), .B1(new_n634), .B2(new_n825), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n840), .B1(new_n639), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n645), .B1(new_n921), .B2(new_n893), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n841), .A2(new_n833), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n723), .B(new_n922), .C1(new_n923), .C2(new_n892), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n733), .B1(new_n924), .B2(new_n847), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n769), .B1(new_n925), .B2(new_n851), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n690), .A2(new_n591), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n491), .A2(KEYINPUT57), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n919), .A2(KEYINPUT57), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n724), .ZN(new_n931));
  INV_X1    g730(.A(new_n885), .ZN(new_n932));
  OAI21_X1  g731(.A(G148gat), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g732(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n906), .A2(new_n724), .A3(new_n908), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n368), .A2(KEYINPUT59), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n919), .A2(new_n932), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n368), .A3(new_n724), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1345gat));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n663), .A3(new_n670), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n906), .A2(new_n670), .A3(new_n908), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n663), .ZN(G1346gat));
  INV_X1    g743(.A(G162gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n939), .A2(new_n945), .A3(new_n733), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n906), .A2(new_n733), .A3(new_n908), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(new_n945), .ZN(G1347gat));
  AOI21_X1  g747(.A(new_n695), .B1(new_n852), .B2(new_n858), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(new_n699), .A3(new_n509), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n723), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n724), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n269), .A3(new_n670), .ZN(new_n955));
  XNOR2_X1  g754(.A(KEYINPUT60), .B(G183gat), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(G1350gat));
  NAND2_X1  g756(.A1(new_n950), .A2(new_n733), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT123), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n235), .B1(new_n959), .B2(KEYINPUT61), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n958), .B(new_n960), .C1(new_n959), .C2(KEYINPUT61), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(G190gat), .B2(new_n958), .ZN(new_n962));
  AOI211_X1 g761(.A(new_n959), .B(KEYINPUT61), .C1(new_n958), .C2(G190gat), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n962), .A2(new_n963), .ZN(G1351gat));
  AND4_X1   g763(.A1(new_n699), .A2(new_n949), .A3(new_n471), .A4(new_n717), .ZN(new_n965));
  INV_X1    g764(.A(G197gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n723), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n695), .A2(new_n492), .A3(new_n323), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n928), .A2(new_n929), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n968), .B(new_n969), .C1(new_n884), .C2(new_n889), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT124), .B1(new_n970), .B2(new_n591), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G197gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n970), .A2(KEYINPUT124), .A3(new_n591), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n976), .B(new_n967), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1352gat));
  INV_X1    g777(.A(new_n931), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n968), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n979), .A2(new_n982), .A3(new_n968), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n981), .A2(G204gat), .A3(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  AOI21_X1  g784(.A(G204gat), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n965), .A2(new_n724), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n984), .A2(new_n989), .ZN(G1353gat));
  OAI21_X1  g789(.A(G211gat), .B1(new_n970), .B2(new_n769), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  NAND3_X1  g791(.A1(new_n965), .A2(new_n339), .A3(new_n670), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1354gat));
  NAND3_X1  g793(.A1(new_n965), .A2(new_n340), .A3(new_n733), .ZN(new_n995));
  OAI21_X1  g794(.A(G218gat), .B1(new_n970), .B2(new_n688), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1355gat));
endmodule


