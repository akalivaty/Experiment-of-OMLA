//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(G230gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT10), .ZN(new_n206));
  AND2_X1   g005(.A1(G71gat), .A2(G78gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  XOR2_X1   g007(.A(G57gat), .B(G64gat), .Z(new_n209));
  AOI211_X1 g008(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(KEYINPUT9), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n207), .B1(KEYINPUT9), .B2(new_n208), .ZN(new_n211));
  INV_X1    g010(.A(G64gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G57gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT88), .B(G57gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G64gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n219), .A2(G85gat), .A3(G92gat), .A4(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n222));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n222), .A2(new_n223), .B1(new_n224), .B2(KEYINPUT8), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n221), .B(new_n225), .C1(G85gat), .C2(G92gat), .ZN(new_n226));
  XOR2_X1   g025(.A(G99gat), .B(G106gat), .Z(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT93), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n229), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT94), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(KEYINPUT94), .A3(new_n231), .A4(new_n232), .ZN(new_n236));
  AOI211_X1 g035(.A(new_n206), .B(new_n218), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n226), .A2(KEYINPUT95), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(new_n227), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n217), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n233), .B2(new_n217), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n205), .B1(new_n237), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G120gat), .B(G148gat), .ZN(new_n245));
  INV_X1    g044(.A(G176gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G204gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n244), .B(new_n250), .C1(new_n205), .C2(new_n241), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n233), .A2(new_n234), .ZN(new_n252));
  INV_X1    g051(.A(new_n236), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT10), .B(new_n217), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n241), .A2(new_n242), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n204), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n241), .A2(new_n205), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n249), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n235), .A2(new_n236), .ZN(new_n263));
  INV_X1    g062(.A(G29gat), .ZN(new_n264));
  INV_X1    g063(.A(G36gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(G29gat), .B2(G36gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT14), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G43gat), .B(G50gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT15), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT81), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G43gat), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(KEYINPUT81), .A3(G50gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT80), .B(KEYINPUT15), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n269), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n271), .B2(new_n269), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT82), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT17), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(KEYINPUT82), .B2(new_n279), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n285), .A2(KEYINPUT17), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(KEYINPUT17), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n263), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n235), .B2(new_n236), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AND4_X1   g094(.A1(new_n262), .A2(new_n292), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n291), .B2(new_n263), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n262), .B1(new_n297), .B2(new_n293), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n261), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n297), .A2(new_n262), .A3(new_n293), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(G218gat), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G134gat), .B(G162gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n299), .A2(new_n303), .A3(new_n304), .A4(new_n308), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT16), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(G1gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G1gat), .B2(new_n313), .ZN(new_n316));
  INV_X1    g115(.A(G8gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT85), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(KEYINPUT85), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n217), .A2(KEYINPUT21), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n217), .A2(KEYINPUT21), .ZN(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n322), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G183gat), .B(G211gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT90), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n326), .B(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT89), .B(G155gat), .Z(new_n332));
  NAND2_X1  g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n331), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n312), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  OAI21_X1  g139(.A(G127gat), .B1(new_n340), .B2(KEYINPUT1), .ZN(new_n341));
  INV_X1    g140(.A(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G113gat), .ZN(new_n343));
  INV_X1    g142(.A(G113gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT1), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n324), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n341), .A2(new_n348), .A3(G134gat), .ZN(new_n349));
  AOI21_X1  g148(.A(G134gat), .B1(new_n341), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n339), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G134gat), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n340), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n324), .B1(new_n346), .B2(new_n347), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n341), .A2(new_n348), .A3(G134gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G155gat), .B(G162gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G141gat), .B(G148gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  AND2_X1   g163(.A1(KEYINPUT72), .A2(G155gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(KEYINPUT72), .A2(G155gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n364), .B1(new_n367), .B2(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n360), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(KEYINPUT72), .A2(G155gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(G162gat), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n369), .A3(KEYINPUT2), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n358), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n363), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n351), .A2(new_n357), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n365), .A2(new_n366), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT73), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n382), .A2(new_n376), .A3(new_n358), .A4(new_n360), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(new_n363), .A3(new_n355), .A4(new_n356), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n363), .C1(new_n370), .C2(new_n377), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n393), .A2(new_n357), .A3(new_n351), .A4(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n387), .B1(new_n384), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n378), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n383), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT66), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n349), .A2(new_n350), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT66), .B1(new_n355), .B2(new_n356), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n392), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  AND4_X1   g208(.A1(new_n392), .A2(new_n408), .A3(new_n398), .A4(new_n396), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G57gat), .ZN(new_n414));
  INV_X1    g213(.A(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n384), .A2(new_n397), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n404), .B1(new_n349), .B2(new_n350), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n355), .A2(KEYINPUT66), .A3(new_n356), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n401), .B2(new_n402), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n396), .B(new_n417), .C1(new_n421), .C2(KEYINPUT4), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n422), .A2(new_n387), .A3(new_n389), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n411), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425));
  INV_X1    g224(.A(new_n416), .ZN(new_n426));
  INV_X1    g225(.A(new_n358), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n368), .B2(new_n369), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n359), .B1(new_n429), .B2(KEYINPUT73), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n400), .B(new_n362), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT75), .B1(new_n383), .B2(new_n363), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n433), .A2(new_n397), .A3(new_n420), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n396), .A2(new_n398), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT76), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n408), .A2(new_n392), .A3(new_n398), .A4(new_n396), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n390), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n387), .A3(new_n389), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n426), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT6), .B(new_n426), .C1(new_n438), .C2(new_n439), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G197gat), .B(G204gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT68), .B(KEYINPUT22), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G211gat), .B(G218gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G211gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n261), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n447), .B(new_n444), .C1(new_n445), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT69), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n449), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458));
  NAND2_X1  g257(.A1(G183gat), .A2(G190gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT64), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT24), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(G183gat), .B2(G190gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G169gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n246), .A3(KEYINPUT23), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT23), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(G169gat), .B2(G176gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n458), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(KEYINPUT25), .C1(new_n464), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n471), .ZN(new_n479));
  NOR3_X1   g278(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT28), .A3(new_n262), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n262), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n481), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n459), .ZN(new_n490));
  NAND2_X1  g289(.A1(G226gat), .A2(G233gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n477), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G183gat), .A2(G190gat), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n494), .B(new_n481), .C1(new_n485), .C2(new_n488), .ZN(new_n495));
  NOR2_X1   g294(.A1(G183gat), .A2(G190gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n494), .B2(KEYINPUT24), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT64), .B1(new_n494), .B2(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n460), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT25), .B1(new_n500), .B2(new_n474), .ZN(new_n501));
  INV_X1    g300(.A(new_n463), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n502), .A2(new_n475), .A3(new_n496), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n503), .A2(new_n472), .A3(new_n458), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT65), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n462), .A2(new_n465), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n472), .B1(new_n507), .B2(new_n497), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n506), .B(new_n476), .C1(new_n508), .C2(KEYINPUT25), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n495), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n492), .A2(KEYINPUT29), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n457), .B(new_n493), .C1(new_n510), .C2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G8gat), .B(G36gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(new_n212), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G92gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n477), .B2(new_n490), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n510), .B2(new_n492), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n513), .B(new_n516), .C1(new_n518), .C2(new_n457), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT30), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n454), .A2(new_n456), .ZN(new_n522));
  AOI211_X1 g321(.A(new_n491), .B(new_n495), .C1(new_n505), .C2(new_n509), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n517), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n513), .ZN(new_n525));
  INV_X1    g324(.A(new_n516), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n519), .A2(KEYINPUT70), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n443), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n506), .B1(new_n473), .B2(new_n476), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT65), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n490), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n407), .ZN(new_n536));
  INV_X1    g335(.A(G227gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(new_n203), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n420), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT32), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G43gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G99gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(KEYINPUT33), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT33), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n540), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT67), .A3(new_n541), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT67), .B1(new_n550), .B2(new_n541), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n539), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n510), .A2(new_n420), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n555), .A2(new_n556), .B1(new_n537), .B2(new_n203), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT34), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n559));
  OAI221_X1 g358(.A(new_n559), .B1(new_n537), .B2(new_n203), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G22gat), .B(G50gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n395), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n457), .ZN(new_n567));
  NAND2_X1  g366(.A1(G228gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n452), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n452), .A2(new_n569), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n449), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT3), .B1(new_n572), .B2(new_n565), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n567), .B(new_n568), .C1(new_n403), .C2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n568), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n522), .B1(new_n565), .B2(new_n395), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT3), .B1(new_n453), .B2(new_n565), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(new_n383), .B2(new_n363), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n574), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n574), .B2(new_n579), .ZN(new_n583));
  XOR2_X1   g382(.A(G78gat), .B(G106gat), .Z(new_n584));
  NOR3_X1   g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n574), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT31), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n588), .B2(new_n581), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n564), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n582), .B2(new_n583), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n581), .A3(new_n586), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n563), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n540), .A2(new_n549), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n541), .A2(new_n595), .A3(new_n545), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n551), .ZN(new_n599));
  INV_X1    g398(.A(new_n561), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n547), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n562), .A2(new_n594), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT35), .B1(new_n532), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n599), .B2(new_n547), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n561), .B(new_n546), .C1(new_n598), .C2(new_n551), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n530), .B1(new_n441), .B2(new_n442), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .A4(new_n594), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n604), .B2(new_n605), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n562), .A2(new_n601), .A3(KEYINPUT36), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n594), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n532), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n513), .B(new_n617), .C1(new_n518), .C2(new_n457), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n524), .A2(KEYINPUT79), .A3(new_n617), .A4(new_n513), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n522), .B(new_n493), .C1(new_n510), .C2(new_n512), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n624), .B(KEYINPUT37), .C1(new_n518), .C2(new_n522), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n622), .A2(new_n623), .A3(new_n526), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n525), .A2(KEYINPUT37), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n526), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n519), .A2(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n441), .A2(new_n442), .A3(new_n626), .A4(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n385), .A2(new_n387), .ZN(new_n634));
  AOI211_X1 g433(.A(new_n633), .B(new_n634), .C1(new_n422), .C2(new_n387), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n422), .A2(new_n633), .A3(new_n387), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n416), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n632), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n422), .A2(new_n387), .ZN(new_n639));
  INV_X1    g438(.A(new_n634), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(KEYINPUT39), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(KEYINPUT40), .A3(new_n416), .A4(new_n636), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n638), .A2(new_n642), .A3(new_n440), .A4(new_n530), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(new_n594), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n614), .A2(new_n616), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n610), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n287), .B1(new_n320), .B2(new_n319), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n291), .B2(new_n318), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT84), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n650), .B(KEYINPUT13), .Z(new_n654));
  AND3_X1   g453(.A1(new_n287), .A2(new_n320), .A3(new_n319), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n654), .B1(new_n655), .B2(new_n647), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT86), .B(new_n654), .C1(new_n655), .C2(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(KEYINPUT18), .A3(new_n650), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n653), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G113gat), .B(G141gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G197gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT11), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n467), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT12), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n653), .A2(new_n660), .A3(new_n667), .A4(new_n661), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n338), .B1(new_n646), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  AOI211_X1 g472(.A(KEYINPUT87), .B(new_n673), .C1(new_n610), .C2(new_n645), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n260), .B(new_n337), .C1(new_n672), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT97), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n643), .A2(new_n594), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n613), .A2(new_n612), .B1(new_n677), .B2(new_n631), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n678), .A2(new_n616), .B1(new_n603), .B2(new_n609), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT87), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n646), .A2(new_n338), .A3(new_n671), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n260), .A4(new_n337), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n443), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n530), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n689), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n314), .A2(new_n317), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n690), .A2(new_n691), .B1(G8gat), .B2(new_n689), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(G1325gat));
  AOI21_X1  g495(.A(G15gat), .B1(new_n685), .B2(new_n606), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n614), .B1(new_n676), .B2(new_n684), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(G15gat), .B2(new_n698), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n615), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT98), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n704), .A3(new_n615), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n685), .B2(new_n615), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT98), .B(new_n594), .C1(new_n676), .C2(new_n684), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT43), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n700), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(new_n701), .A3(new_n705), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n707), .B2(new_n708), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n712), .A3(G22gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(G1327gat));
  NOR2_X1   g513(.A1(new_n335), .A2(new_n259), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n312), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n680), .B2(new_n681), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n264), .A3(new_n686), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n310), .A2(new_n311), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n679), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n720), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n671), .B(new_n715), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G29gat), .B1(new_n725), .B2(new_n443), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n726), .ZN(G1328gat));
  INV_X1    g526(.A(new_n725), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n265), .B1(new_n728), .B2(new_n530), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n265), .A3(new_n530), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT99), .B1(new_n730), .B2(KEYINPUT46), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(KEYINPUT99), .A3(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n732), .B(new_n733), .C1(KEYINPUT46), .C2(new_n730), .ZN(G1329gat));
  OAI21_X1  g533(.A(G43gat), .B1(new_n725), .B2(new_n614), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n604), .A2(new_n605), .A3(G43gat), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT100), .B1(new_n717), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n717), .A2(KEYINPUT100), .A3(new_n736), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(KEYINPUT47), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT101), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n739), .B2(new_n737), .ZN(new_n742));
  INV_X1    g541(.A(new_n737), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(KEYINPUT101), .A3(new_n738), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n744), .A3(new_n735), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n745), .A2(KEYINPUT102), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT102), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n615), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n725), .B2(new_n594), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(G50gat), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n717), .A2(new_n754), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n755), .A2(KEYINPUT104), .A3(new_n594), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT104), .B1(new_n755), .B2(new_n594), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n753), .A2(new_n756), .A3(new_n757), .A4(KEYINPUT48), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT103), .B(KEYINPUT48), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n754), .B1(new_n728), .B2(new_n615), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n755), .A2(new_n594), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n762), .ZN(G1331gat));
  AND4_X1   g562(.A1(new_n259), .A2(new_n646), .A3(new_n673), .A4(new_n337), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n686), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(new_n214), .Z(G1332gat));
  AOI21_X1  g565(.A(new_n531), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT106), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT107), .Z(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1333gat));
  INV_X1    g571(.A(new_n614), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n764), .A2(G71gat), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n764), .A2(new_n606), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(G71gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT108), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g577(.A1(new_n764), .A2(new_n615), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n671), .A2(new_n335), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT109), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n721), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n259), .ZN(new_n786));
  AOI21_X1  g585(.A(G85gat), .B1(new_n786), .B2(new_n686), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n259), .B(new_n782), .C1(new_n723), .C2(new_n724), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(new_n415), .A3(new_n443), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n787), .A2(KEYINPUT110), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n787), .B2(new_n789), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1336gat));
  NOR3_X1   g591(.A1(new_n260), .A2(G92gat), .A3(new_n531), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G92gat), .B1(new_n788), .B2(new_n531), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n784), .A2(KEYINPUT111), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n783), .B(new_n799), .Z(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n798), .B1(new_n801), .B2(new_n795), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT112), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n797), .B2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1337gat));
  NOR3_X1   g606(.A1(new_n788), .A2(new_n544), .A3(new_n614), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n606), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n544), .ZN(G1338gat));
  NOR2_X1   g609(.A1(new_n594), .A2(G106gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n785), .A2(new_n259), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT113), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(G106gat), .B1(new_n788), .B2(new_n594), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n259), .A3(new_n811), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n815), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n814), .B2(new_n818), .ZN(G1339gat));
  OR2_X1    g618(.A1(new_n655), .A2(new_n647), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n648), .A2(new_n650), .B1(new_n820), .B2(new_n654), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n666), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n259), .A2(new_n670), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n254), .A2(new_n204), .A3(new_n255), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n244), .A2(KEYINPUT54), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n250), .B1(new_n256), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT55), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n251), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n823), .B1(new_n673), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n720), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n670), .A2(new_n822), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n310), .B2(new_n311), .ZN(new_n836));
  INV_X1    g635(.A(new_n832), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n335), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NOR4_X1   g638(.A1(new_n312), .A2(new_n336), .A3(new_n259), .A4(new_n671), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n686), .A2(new_n531), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n602), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n673), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n344), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n845), .A2(new_n260), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n342), .ZN(G1341gat));
  NOR3_X1   g648(.A1(new_n845), .A2(new_n324), .A3(new_n336), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT114), .ZN(new_n851));
  INV_X1    g650(.A(new_n845), .ZN(new_n852));
  AOI21_X1  g651(.A(G127gat), .B1(new_n852), .B2(new_n335), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(G1342gat));
  NAND2_X1  g653(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n312), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT115), .Z(new_n858));
  XNOR2_X1  g657(.A(new_n856), .B(new_n858), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n594), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n773), .A2(new_n842), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n864));
  NAND2_X1  g663(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n866));
  OR2_X1    g665(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n251), .A3(new_n671), .A4(new_n831), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n312), .B1(new_n869), .B2(new_n823), .ZN(new_n870));
  INV_X1    g669(.A(new_n838), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n336), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n840), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n594), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n862), .B(new_n863), .C1(new_n861), .C2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n875), .B2(new_n673), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n843), .A2(new_n615), .A3(new_n614), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n673), .A2(G141gat), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT118), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT58), .ZN(G1344gat));
  OR3_X1    g681(.A1(new_n877), .A2(G148gat), .A3(new_n260), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n884), .B(G148gat), .C1(new_n875), .C2(new_n260), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(KEYINPUT57), .B2(new_n874), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n259), .A3(new_n863), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n886), .B2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(new_n367), .B1(new_n875), .B2(new_n336), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n877), .A2(new_n367), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n336), .B2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n875), .B2(new_n720), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n380), .A3(new_n312), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n686), .A2(new_n531), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n844), .B(new_n898), .C1(new_n839), .C2(new_n840), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n720), .A2(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n873), .B1(new_n901), .B2(new_n335), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n844), .A4(new_n898), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n467), .B1(new_n905), .B2(new_n671), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT120), .ZN(new_n907));
  INV_X1    g706(.A(new_n899), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n467), .A3(new_n671), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1348gat));
  INV_X1    g709(.A(new_n905), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n246), .A3(new_n260), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n246), .B1(new_n899), .B2(new_n260), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT121), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n912), .A2(new_n914), .ZN(G1349gat));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(new_n905), .B2(new_n335), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918));
  AOI211_X1 g717(.A(new_n918), .B(new_n336), .C1(new_n900), .C2(new_n904), .ZN(new_n919));
  INV_X1    g718(.A(G183gat), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n908), .A2(new_n484), .A3(new_n335), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT123), .B(new_n916), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n917), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n335), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(G183gat), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n916), .A2(KEYINPUT123), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n916), .A2(KEYINPUT123), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .A4(new_n922), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n924), .A2(new_n930), .ZN(G1350gat));
  AOI21_X1  g730(.A(new_n262), .B1(new_n905), .B2(new_n312), .ZN(new_n932));
  XNOR2_X1  g731(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n908), .A2(new_n262), .A3(new_n312), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1351gat));
  NAND2_X1  g735(.A1(new_n614), .A2(new_n898), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n888), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n673), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n860), .A2(new_n938), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n673), .A2(G197gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  AND2_X1   g742(.A1(new_n888), .A2(new_n259), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n248), .B1(new_n944), .B2(new_n938), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n860), .A2(new_n248), .A3(new_n938), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n260), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n946), .B(KEYINPUT62), .C1(new_n948), .C2(new_n260), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT126), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n888), .A2(new_n259), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n955), .B2(new_n937), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n956), .A2(new_n957), .A3(new_n951), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n958), .ZN(G1353gat));
  NAND4_X1  g758(.A1(new_n860), .A2(new_n450), .A3(new_n335), .A4(new_n938), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n888), .A2(new_n335), .A3(new_n938), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  OAI21_X1  g763(.A(new_n261), .B1(new_n941), .B2(new_n720), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n939), .A2(new_n261), .A3(new_n720), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(G1355gat));
endmodule


