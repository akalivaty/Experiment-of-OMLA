

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U321 ( .A(n307), .B(n306), .ZN(n522) );
  XOR2_X1 U322 ( .A(n450), .B(KEYINPUT41), .Z(n549) );
  XNOR2_X1 U323 ( .A(n296), .B(KEYINPUT89), .ZN(n297) );
  NOR2_X1 U324 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U325 ( .A(n298), .B(n297), .ZN(n423) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n529) );
  INV_X1 U327 ( .A(n529), .ZN(n530) );
  XNOR2_X1 U328 ( .A(n454), .B(G218GAT), .ZN(n455) );
  XNOR2_X1 U329 ( .A(n451), .B(G204GAT), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n480), .B(G43GAT), .ZN(n481) );
  XNOR2_X1 U331 ( .A(n456), .B(n455), .ZN(G1355GAT) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(G1353GAT) );
  XNOR2_X1 U333 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n294) );
  XNOR2_X1 U335 ( .A(G36GAT), .B(KEYINPUT76), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n289), .B(G190GAT), .ZN(n313) );
  XOR2_X1 U337 ( .A(G204GAT), .B(KEYINPUT71), .Z(n291) );
  XNOR2_X1 U338 ( .A(G92GAT), .B(G176GAT), .ZN(n290) );
  XNOR2_X1 U339 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U340 ( .A(G64GAT), .B(n292), .Z(n332) );
  XNOR2_X1 U341 ( .A(n313), .B(n332), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n302) );
  XNOR2_X1 U343 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n295), .B(KEYINPUT88), .ZN(n298) );
  XNOR2_X1 U345 ( .A(G218GAT), .B(G211GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n423), .B(KEYINPUT93), .ZN(n300) );
  NAND2_X1 U347 ( .A1(G226GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U349 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U350 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT17), .B(G169GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(G183GAT), .B(n305), .Z(n443) );
  XNOR2_X1 U354 ( .A(G8GAT), .B(n443), .ZN(n306) );
  XOR2_X1 U355 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n309) );
  XNOR2_X1 U356 ( .A(G92GAT), .B(KEYINPUT75), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(n310), .B(G106GAT), .Z(n312) );
  XOR2_X1 U359 ( .A(G162GAT), .B(G50GAT), .Z(n420) );
  XNOR2_X1 U360 ( .A(n420), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n312), .B(n311), .ZN(n317) );
  XOR2_X1 U362 ( .A(G85GAT), .B(G99GAT), .Z(n333) );
  XOR2_X1 U363 ( .A(n333), .B(n313), .Z(n315) );
  NAND2_X1 U364 ( .A1(G232GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U366 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U367 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n319) );
  XNOR2_X1 U368 ( .A(KEYINPUT67), .B(G43GAT), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U370 ( .A(G29GAT), .B(n320), .Z(n355) );
  XOR2_X1 U371 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n322) );
  XNOR2_X1 U372 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n355), .B(n323), .ZN(n324) );
  XOR2_X1 U375 ( .A(n325), .B(n324), .Z(n575) );
  INV_X1 U376 ( .A(n575), .ZN(n483) );
  XOR2_X1 U377 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n357) );
  XOR2_X1 U378 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .Z(n361) );
  XOR2_X1 U380 ( .A(n428), .B(n361), .Z(n327) );
  NAND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U383 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n329) );
  XNOR2_X1 U384 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U386 ( .A(n331), .B(n330), .Z(n335) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n337) );
  INV_X1 U389 ( .A(KEYINPUT32), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT70), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U392 ( .A(G148GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n415) );
  XOR2_X1 U394 ( .A(n415), .B(KEYINPUT31), .Z(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n450) );
  XOR2_X1 U396 ( .A(G197GAT), .B(G50GAT), .Z(n343) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(G36GAT), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U399 ( .A(KEYINPUT29), .B(G169GAT), .Z(n345) );
  XNOR2_X1 U400 ( .A(G113GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n353) );
  XOR2_X1 U403 ( .A(KEYINPUT68), .B(G8GAT), .Z(n349) );
  XNOR2_X1 U404 ( .A(G1GAT), .B(G22GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U406 ( .A(n364), .B(KEYINPUT30), .Z(n351) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n355), .B(n354), .Z(n505) );
  INV_X1 U411 ( .A(n505), .ZN(n564) );
  NAND2_X1 U412 ( .A1(n549), .A2(n564), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n377) );
  XOR2_X1 U414 ( .A(G64GAT), .B(G183GAT), .Z(n359) );
  XNOR2_X1 U415 ( .A(G78GAT), .B(G71GAT), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U417 ( .A(n360), .B(G211GAT), .Z(n363) );
  XNOR2_X1 U418 ( .A(G155GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U420 ( .A(G127GAT), .B(G15GAT), .Z(n437) );
  XOR2_X1 U421 ( .A(n364), .B(n437), .Z(n366) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n376) );
  XOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n370) );
  XNOR2_X1 U426 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n372) );
  XNOR2_X1 U429 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U432 ( .A(n376), .B(n375), .Z(n580) );
  NOR2_X1 U433 ( .A1(n377), .A2(n580), .ZN(n378) );
  NAND2_X1 U434 ( .A1(n483), .A2(n378), .ZN(n379) );
  XNOR2_X1 U435 ( .A(KEYINPUT47), .B(n379), .ZN(n385) );
  XOR2_X1 U436 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT36), .B(n575), .ZN(n471) );
  NAND2_X1 U438 ( .A1(n471), .A2(n580), .ZN(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n383) );
  INV_X1 U440 ( .A(n450), .ZN(n477) );
  NAND2_X1 U441 ( .A1(n505), .A2(n477), .ZN(n382) );
  NOR2_X1 U442 ( .A1(n383), .A2(n382), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n385), .A2(n384), .ZN(n388) );
  XNOR2_X1 U444 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n386), .B(KEYINPUT114), .ZN(n387) );
  NOR2_X1 U446 ( .A1(n522), .A2(n529), .ZN(n390) );
  XNOR2_X1 U447 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n411) );
  XOR2_X1 U449 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n392) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n410) );
  XOR2_X1 U452 ( .A(G127GAT), .B(G120GAT), .Z(n394) );
  XNOR2_X1 U453 ( .A(G162GAT), .B(G148GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U455 ( .A(G29GAT), .B(G85GAT), .Z(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n406) );
  XOR2_X1 U457 ( .A(G141GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n416) );
  XOR2_X1 U460 ( .A(G113GAT), .B(KEYINPUT83), .Z(n400) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n429) );
  XNOR2_X1 U463 ( .A(n416), .B(n429), .ZN(n404) );
  XOR2_X1 U464 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n402) );
  XNOR2_X1 U465 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n408) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U471 ( .A(n410), .B(n409), .Z(n518) );
  NAND2_X1 U472 ( .A1(n411), .A2(n518), .ZN(n559) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n413) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U476 ( .A(n414), .B(KEYINPUT23), .Z(n418) );
  XNOR2_X1 U477 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n419), .B(G204GAT), .Z(n422) );
  XNOR2_X1 U480 ( .A(n420), .B(G22GAT), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n425) );
  INV_X1 U482 ( .A(n423), .ZN(n424) );
  XOR2_X1 U483 ( .A(n425), .B(n424), .Z(n558) );
  XOR2_X1 U484 ( .A(G176GAT), .B(KEYINPUT65), .Z(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n441) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n435) );
  XNOR2_X1 U492 ( .A(G190GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U494 ( .A(n436), .B(KEYINPUT84), .Z(n439) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X2 U498 ( .A(n443), .B(n442), .Z(n563) );
  INV_X1 U499 ( .A(n563), .ZN(n533) );
  NOR2_X1 U500 ( .A1(n558), .A2(n533), .ZN(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n545) );
  NOR2_X1 U503 ( .A1(n559), .A2(n545), .ZN(n446) );
  XOR2_X1 U504 ( .A(KEYINPUT125), .B(n446), .Z(n579) );
  NAND2_X1 U505 ( .A1(n579), .A2(n564), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n447) );
  XNOR2_X1 U507 ( .A(n447), .B(G197GAT), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(G1352GAT) );
  NAND2_X1 U509 ( .A1(n579), .A2(n450), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n451) );
  NAND2_X1 U511 ( .A1(n579), .A2(n471), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n454) );
  INV_X1 U513 ( .A(KEYINPUT38), .ZN(n479) );
  XNOR2_X1 U514 ( .A(n522), .B(KEYINPUT95), .ZN(n457) );
  XOR2_X1 U515 ( .A(n457), .B(KEYINPUT27), .Z(n466) );
  OR2_X1 U516 ( .A1(n545), .A2(n466), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n563), .A2(n522), .ZN(n458) );
  XNOR2_X1 U518 ( .A(KEYINPUT97), .B(n458), .ZN(n459) );
  NAND2_X1 U519 ( .A1(n459), .A2(n558), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT98), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NAND2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n518), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n465), .B(KEYINPUT99), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n518), .A2(n466), .ZN(n531) );
  NAND2_X1 U526 ( .A1(n563), .A2(n531), .ZN(n467) );
  XOR2_X1 U527 ( .A(KEYINPUT28), .B(n558), .Z(n496) );
  NOR2_X1 U528 ( .A1(n467), .A2(n496), .ZN(n468) );
  XOR2_X1 U529 ( .A(KEYINPUT100), .B(n470), .Z(n487) );
  INV_X1 U530 ( .A(n580), .ZN(n472) );
  AND2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n473) );
  AND2_X1 U532 ( .A1(n487), .A2(n473), .ZN(n476) );
  XOR2_X1 U533 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT37), .B(n474), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n517) );
  NAND2_X1 U536 ( .A1(n477), .A2(n564), .ZN(n488) );
  NOR2_X1 U537 ( .A1(n517), .A2(n488), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n503) );
  NOR2_X1 U539 ( .A1(n563), .A2(n503), .ZN(n482) );
  INV_X1 U540 ( .A(KEYINPUT40), .ZN(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n485) );
  NAND2_X1 U542 ( .A1(n483), .A2(n580), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U544 ( .A1(n487), .A2(n486), .ZN(n506) );
  NOR2_X1 U545 ( .A1(n506), .A2(n488), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT101), .ZN(n497) );
  NOR2_X1 U547 ( .A1(n518), .A2(n497), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n492), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n522), .A2(n497), .ZN(n493) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n563), .A2(n497), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  INV_X1 U556 ( .A(n496), .ZN(n532) );
  NOR2_X1 U557 ( .A1(n532), .A2(n497), .ZN(n499) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(G1327GAT) );
  NOR2_X1 U560 ( .A1(n503), .A2(n518), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n522), .ZN(n502) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U565 ( .A1(n503), .A2(n532), .ZN(n504) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XNOR2_X1 U567 ( .A(KEYINPUT106), .B(n549), .ZN(n571) );
  NAND2_X1 U568 ( .A1(n505), .A2(n571), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n506), .A2(n516), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT107), .B(n507), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n518), .A2(n513), .ZN(n508) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n513), .ZN(n510) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n563), .A2(n513), .ZN(n511) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(n511), .Z(n512) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n532), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  OR2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n518), .A2(n526), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n526), .ZN(n524) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1337GAT) );
  NOR2_X1 U590 ( .A1(n563), .A2(n526), .ZN(n525) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n525), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n532), .A2(n526), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U597 ( .A1(n544), .A2(n534), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n564), .A2(n541), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n571), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n580), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n575), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT117), .Z(n548) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT116), .B(n546), .ZN(n555) );
  NAND2_X1 U613 ( .A1(n555), .A2(n564), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U617 ( .A1(n555), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n580), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT119), .Z(n557) );
  NAND2_X1 U623 ( .A1(n555), .A2(n575), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n566) );
  INV_X1 U626 ( .A(n558), .ZN(n560) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT55), .ZN(n562) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n576), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n569) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(n570), .Z(n573) );
  NAND2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n580), .A2(n576), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1351GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
endmodule

