

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748;

  NAND2_X1 U372 ( .A1(n351), .A2(n404), .ZN(n407) );
  NAND2_X1 U373 ( .A1(n406), .A2(n405), .ZN(n351) );
  XNOR2_X1 U374 ( .A(n369), .B(n499), .ZN(n533) );
  OR2_X1 U375 ( .A1(n392), .A2(n388), .ZN(n538) );
  AND2_X4 U376 ( .A1(n407), .A2(n439), .ZN(n708) );
  NOR2_X2 U377 ( .A1(n681), .A2(n497), .ZN(n406) );
  XNOR2_X2 U378 ( .A(n435), .B(KEYINPUT107), .ZN(n742) );
  XNOR2_X2 U379 ( .A(n729), .B(G146), .ZN(n484) );
  NOR2_X1 U380 ( .A1(n620), .A2(G902), .ZN(n486) );
  XNOR2_X1 U381 ( .A(n434), .B(n433), .ZN(n741) );
  NOR2_X1 U382 ( .A1(n551), .A2(n572), .ZN(n500) );
  NAND2_X1 U383 ( .A1(n372), .A2(n371), .ZN(n592) );
  NOR2_X1 U384 ( .A1(n551), .A2(n649), .ZN(n553) );
  AND2_X1 U385 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U386 ( .A1(n429), .A2(n428), .ZN(n427) );
  XNOR2_X1 U387 ( .A(n459), .B(n458), .ZN(n658) );
  XNOR2_X1 U388 ( .A(n691), .B(n366), .ZN(n692) );
  NAND2_X1 U389 ( .A1(n619), .A2(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U390 ( .A(n478), .B(n437), .ZN(n494) );
  XNOR2_X1 U391 ( .A(G119), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U392 ( .A(n438), .B(G116), .ZN(n437) );
  INV_X1 U393 ( .A(G113), .ZN(n438) );
  XNOR2_X1 U394 ( .A(n487), .B(n398), .ZN(n397) );
  NAND2_X1 U395 ( .A1(n697), .A2(n470), .ZN(n394) );
  XNOR2_X1 U396 ( .A(n589), .B(KEYINPUT22), .ZN(n602) );
  XNOR2_X1 U397 ( .A(n353), .B(n464), .ZN(n714) );
  XNOR2_X1 U398 ( .A(n714), .B(n465), .ZN(n490) );
  INV_X1 U399 ( .A(KEYINPUT73), .ZN(n465) );
  NAND2_X1 U400 ( .A1(n408), .A2(n722), .ZN(n439) );
  NOR2_X1 U401 ( .A1(n618), .A2(n617), .ZN(n408) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n510) );
  XNOR2_X1 U403 ( .A(n460), .B(KEYINPUT4), .ZN(n420) );
  INV_X1 U404 ( .A(KEYINPUT66), .ZN(n460) );
  XNOR2_X1 U405 ( .A(n426), .B(G125), .ZN(n489) );
  INV_X1 U406 ( .A(G146), .ZN(n426) );
  INV_X1 U407 ( .A(n741), .ZN(n379) );
  NOR2_X1 U408 ( .A1(n741), .A2(KEYINPUT44), .ZN(n381) );
  XOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n493) );
  XNOR2_X1 U410 ( .A(n491), .B(n489), .ZN(n417) );
  NAND2_X1 U411 ( .A1(n377), .A2(n354), .ZN(n376) );
  INV_X1 U412 ( .A(n430), .ZN(n377) );
  NAND2_X1 U413 ( .A1(n374), .A2(n354), .ZN(n373) );
  NAND2_X1 U414 ( .A1(n427), .A2(n375), .ZN(n374) );
  INV_X1 U415 ( .A(n584), .ZN(n375) );
  XNOR2_X1 U416 ( .A(n401), .B(G478), .ZN(n555) );
  OR2_X1 U417 ( .A1(n706), .A2(G902), .ZN(n401) );
  INV_X1 U418 ( .A(G902), .ZN(n390) );
  XNOR2_X1 U419 ( .A(n538), .B(KEYINPUT1), .ZN(n576) );
  XNOR2_X1 U420 ( .A(n484), .B(n485), .ZN(n620) );
  XNOR2_X1 U421 ( .A(n483), .B(n368), .ZN(n485) );
  XNOR2_X1 U422 ( .A(n494), .B(n482), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n494), .B(n436), .ZN(n713) );
  XNOR2_X1 U424 ( .A(G122), .B(KEYINPUT16), .ZN(n436) );
  INV_X1 U425 ( .A(KEYINPUT39), .ZN(n552) );
  XNOR2_X1 U426 ( .A(n457), .B(n456), .ZN(n458) );
  NOR2_X1 U427 ( .A1(n602), .A2(n590), .ZN(n608) );
  XNOR2_X1 U428 ( .A(n484), .B(n440), .ZN(n697) );
  XNOR2_X1 U429 ( .A(n466), .B(n469), .ZN(n440) );
  INV_X1 U430 ( .A(n490), .ZN(n466) );
  NOR2_X1 U431 ( .A1(n736), .A2(G952), .ZN(n712) );
  INV_X1 U432 ( .A(n684), .ZN(n378) );
  INV_X1 U433 ( .A(n742), .ZN(n382) );
  NAND2_X1 U434 ( .A1(n416), .A2(n415), .ZN(n414) );
  INV_X1 U435 ( .A(n529), .ZN(n415) );
  NAND2_X1 U436 ( .A1(n662), .A2(n569), .ZN(n487) );
  INV_X1 U437 ( .A(KEYINPUT30), .ZN(n398) );
  XOR2_X1 U438 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n480) );
  XNOR2_X1 U439 ( .A(G131), .B(G101), .ZN(n482) );
  XNOR2_X1 U440 ( .A(n489), .B(n425), .ZN(n503) );
  INV_X1 U441 ( .A(KEYINPUT10), .ZN(n425) );
  XOR2_X1 U442 ( .A(G104), .B(G122), .Z(n512) );
  XNOR2_X1 U443 ( .A(n491), .B(n463), .ZN(n729) );
  XNOR2_X1 U444 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U445 ( .A(G137), .B(KEYINPUT70), .Z(n462) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n471) );
  AND2_X1 U447 ( .A1(n658), .A2(n422), .ZN(n541) );
  NOR2_X1 U448 ( .A1(n659), .A2(n529), .ZN(n422) );
  XNOR2_X1 U449 ( .A(G119), .B(G137), .ZN(n449) );
  XOR2_X1 U450 ( .A(KEYINPUT23), .B(G110), .Z(n450) );
  XNOR2_X1 U451 ( .A(n503), .B(n423), .ZN(n446) );
  XNOR2_X1 U452 ( .A(n444), .B(n424), .ZN(n423) );
  INV_X1 U453 ( .A(KEYINPUT94), .ZN(n424) );
  XNOR2_X1 U454 ( .A(KEYINPUT95), .B(KEYINPUT24), .ZN(n444) );
  XNOR2_X1 U455 ( .A(n520), .B(G107), .ZN(n403) );
  XOR2_X1 U456 ( .A(KEYINPUT7), .B(G122), .Z(n520) );
  XNOR2_X1 U457 ( .A(n370), .B(n496), .ZN(n691) );
  XNOR2_X1 U458 ( .A(n417), .B(n490), .ZN(n370) );
  XNOR2_X1 U459 ( .A(n386), .B(n364), .ZN(n610) );
  NAND2_X1 U460 ( .A1(n352), .A2(n430), .ZN(n371) );
  AND2_X1 U461 ( .A1(n376), .A2(n373), .ZN(n372) );
  NOR2_X1 U462 ( .A1(n664), .A2(n602), .ZN(n603) );
  NAND2_X1 U463 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U464 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U465 ( .A(n604), .ZN(n662) );
  XNOR2_X1 U466 ( .A(n699), .B(n367), .ZN(n700) );
  XNOR2_X1 U467 ( .A(n554), .B(KEYINPUT40), .ZN(n746) );
  XNOR2_X1 U468 ( .A(n609), .B(KEYINPUT32), .ZN(n433) );
  NAND2_X1 U469 ( .A1(n608), .A2(n607), .ZN(n434) );
  INV_X1 U470 ( .A(KEYINPUT78), .ZN(n609) );
  INV_X1 U471 ( .A(KEYINPUT109), .ZN(n412) );
  AND2_X1 U472 ( .A1(n418), .A2(n359), .ZN(n625) );
  XNOR2_X1 U473 ( .A(n608), .B(KEYINPUT86), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n695), .B(n400), .ZN(n698) );
  XNOR2_X1 U475 ( .A(n697), .B(n696), .ZN(n400) );
  NOR2_X1 U476 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U477 ( .A1(n419), .A2(n356), .ZN(n681) );
  AND2_X1 U478 ( .A1(n427), .A2(n361), .ZN(n352) );
  XOR2_X1 U479 ( .A(G107), .B(G104), .Z(n353) );
  XOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT0), .Z(n354) );
  AND2_X1 U481 ( .A1(n556), .A2(n555), .ZN(n355) );
  AND2_X1 U482 ( .A1(n743), .A2(n645), .ZN(n356) );
  AND2_X1 U483 ( .A1(n384), .A2(n383), .ZN(n357) );
  AND2_X1 U484 ( .A1(n382), .A2(n379), .ZN(n358) );
  AND2_X1 U485 ( .A1(n605), .A2(n606), .ZN(n359) );
  AND2_X1 U486 ( .A1(n658), .A2(n604), .ZN(n360) );
  NOR2_X1 U487 ( .A1(n584), .A2(n354), .ZN(n361) );
  NOR2_X1 U488 ( .A1(n405), .A2(n378), .ZN(n362) );
  XOR2_X1 U489 ( .A(KEYINPUT75), .B(KEYINPUT34), .Z(n363) );
  XOR2_X1 U490 ( .A(KEYINPUT35), .B(KEYINPUT85), .Z(n364) );
  XOR2_X1 U491 ( .A(n620), .B(KEYINPUT62), .Z(n365) );
  XNOR2_X1 U492 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n366) );
  XNOR2_X1 U493 ( .A(KEYINPUT59), .B(KEYINPUT91), .ZN(n367) );
  NAND2_X1 U494 ( .A1(n691), .A2(n497), .ZN(n369) );
  NAND2_X1 U495 ( .A1(n430), .A2(n427), .ZN(n583) );
  NAND2_X1 U496 ( .A1(n592), .A2(n588), .ZN(n589) );
  XNOR2_X1 U497 ( .A(n615), .B(KEYINPUT45), .ZN(n405) );
  NAND2_X1 U498 ( .A1(n357), .A2(n380), .ZN(n612) );
  NAND2_X1 U499 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U500 ( .A1(n741), .A2(KEYINPUT44), .ZN(n383) );
  NAND2_X1 U501 ( .A1(n742), .A2(KEYINPUT44), .ZN(n384) );
  NAND2_X1 U502 ( .A1(n358), .A2(n740), .ZN(n611) );
  XNOR2_X2 U503 ( .A(n385), .B(n420), .ZN(n491) );
  XNOR2_X1 U504 ( .A(n385), .B(n403), .ZN(n521) );
  XNOR2_X2 U505 ( .A(n421), .B(G143), .ZN(n385) );
  NAND2_X1 U506 ( .A1(n610), .A2(KEYINPUT44), .ZN(n586) );
  NAND2_X1 U507 ( .A1(n387), .A2(n355), .ZN(n386) );
  XNOR2_X1 U508 ( .A(n585), .B(n363), .ZN(n387) );
  NOR2_X1 U509 ( .A1(n697), .A2(n389), .ZN(n388) );
  INV_X1 U510 ( .A(n470), .ZN(n391) );
  NAND2_X1 U511 ( .A1(n470), .A2(G902), .ZN(n393) );
  NOR2_X2 U512 ( .A1(n702), .A2(n712), .ZN(n704) );
  XNOR2_X1 U513 ( .A(n395), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U514 ( .A1(n694), .A2(n712), .ZN(n395) );
  XNOR2_X2 U515 ( .A(n396), .B(n567), .ZN(n419) );
  NAND2_X1 U516 ( .A1(n565), .A2(n566), .ZN(n396) );
  NAND2_X1 U517 ( .A1(n745), .A2(n746), .ZN(n563) );
  NAND2_X1 U518 ( .A1(n488), .A2(n397), .ZN(n551) );
  NAND2_X1 U519 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U520 ( .A1(n402), .A2(n360), .ZN(n435) );
  XNOR2_X1 U521 ( .A(n603), .B(KEYINPUT106), .ZN(n402) );
  NOR2_X1 U522 ( .A1(n647), .A2(n659), .ZN(n588) );
  XNOR2_X1 U523 ( .A(n557), .B(KEYINPUT105), .ZN(n647) );
  INV_X1 U524 ( .A(KEYINPUT64), .ZN(n409) );
  XNOR2_X2 U525 ( .A(n409), .B(G953), .ZN(n736) );
  NAND2_X1 U526 ( .A1(n736), .A2(G234), .ZN(n448) );
  NAND2_X1 U527 ( .A1(n748), .A2(n527), .ZN(n528) );
  XNOR2_X2 U528 ( .A(n410), .B(KEYINPUT110), .ZN(n748) );
  NAND2_X1 U529 ( .A1(n411), .A2(n355), .ZN(n410) );
  XNOR2_X1 U530 ( .A(n500), .B(n412), .ZN(n411) );
  NOR2_X1 U531 ( .A1(n658), .A2(n414), .ZN(n413) );
  AND2_X1 U532 ( .A1(n538), .A2(n413), .ZN(n477) );
  INV_X1 U533 ( .A(n659), .ZN(n416) );
  NAND2_X1 U534 ( .A1(n665), .A2(n538), .ZN(n595) );
  NOR2_X1 U535 ( .A1(n658), .A2(n659), .ZN(n665) );
  NAND2_X1 U536 ( .A1(n419), .A2(n743), .ZN(n618) );
  XNOR2_X2 U537 ( .A(G128), .B(KEYINPUT79), .ZN(n421) );
  NOR2_X1 U538 ( .A1(n591), .A2(n587), .ZN(n578) );
  XNOR2_X2 U539 ( .A(n486), .B(G472), .ZN(n604) );
  INV_X1 U540 ( .A(n658), .ZN(n606) );
  NAND2_X1 U541 ( .A1(n662), .A2(n541), .ZN(n531) );
  NAND2_X1 U542 ( .A1(n533), .A2(n535), .ZN(n432) );
  NAND2_X1 U543 ( .A1(n429), .A2(n569), .ZN(n542) );
  NOR2_X1 U544 ( .A1(n653), .A2(n535), .ZN(n428) );
  INV_X1 U545 ( .A(n533), .ZN(n429) );
  NAND2_X1 U546 ( .A1(n653), .A2(n535), .ZN(n431) );
  NAND2_X1 U547 ( .A1(n683), .A2(n439), .ZN(n685) );
  NAND2_X1 U548 ( .A1(n576), .A2(n665), .ZN(n591) );
  XNOR2_X1 U549 ( .A(n621), .B(n365), .ZN(n623) );
  INV_X1 U550 ( .A(KEYINPUT71), .ZN(n549) );
  INV_X1 U551 ( .A(KEYINPUT48), .ZN(n567) );
  INV_X1 U552 ( .A(G134), .ZN(n461) );
  XNOR2_X1 U553 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U554 ( .A(n712), .ZN(n622) );
  NAND2_X1 U555 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U556 ( .A(G902), .B(KEYINPUT15), .Z(n619) );
  INV_X1 U557 ( .A(n619), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(G234), .ZN(n442) );
  XNOR2_X1 U559 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U560 ( .A(n442), .B(n441), .ZN(n455) );
  NAND2_X1 U561 ( .A1(n455), .A2(G221), .ZN(n443) );
  XNOR2_X1 U562 ( .A(n443), .B(KEYINPUT21), .ZN(n659) );
  XNOR2_X1 U563 ( .A(G128), .B(G140), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n446), .B(n445), .ZN(n454) );
  XNOR2_X1 U565 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n447) );
  XNOR2_X1 U566 ( .A(n448), .B(n447), .ZN(n523) );
  AND2_X1 U567 ( .A1(G221), .A2(n523), .ZN(n452) );
  XNOR2_X1 U568 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n454), .B(n453), .ZN(n710) );
  NOR2_X1 U570 ( .A1(G902), .A2(n710), .ZN(n459) );
  NAND2_X1 U571 ( .A1(G217), .A2(n455), .ZN(n457) );
  XNOR2_X1 U572 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n456) );
  XNOR2_X1 U573 ( .A(G101), .B(G110), .ZN(n464) );
  XOR2_X1 U574 ( .A(G131), .B(G140), .Z(n501) );
  XOR2_X1 U575 ( .A(n501), .B(KEYINPUT93), .Z(n468) );
  NAND2_X1 U576 ( .A1(G227), .A2(n736), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U578 ( .A(KEYINPUT72), .B(G469), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U580 ( .A1(G952), .A2(n472), .ZN(n680) );
  NOR2_X1 U581 ( .A1(G953), .A2(n680), .ZN(n582) );
  INV_X1 U582 ( .A(n736), .ZN(n473) );
  AND2_X1 U583 ( .A1(G902), .A2(n472), .ZN(n579) );
  NAND2_X1 U584 ( .A1(n473), .A2(n579), .ZN(n474) );
  NOR2_X1 U585 ( .A1(G900), .A2(n474), .ZN(n475) );
  NOR2_X1 U586 ( .A1(n582), .A2(n475), .ZN(n476) );
  XNOR2_X1 U587 ( .A(KEYINPUT80), .B(n476), .ZN(n529) );
  XNOR2_X1 U588 ( .A(n477), .B(KEYINPUT76), .ZN(n488) );
  NAND2_X1 U589 ( .A1(n510), .A2(G210), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U591 ( .A(n481), .B(KEYINPUT5), .Z(n483) );
  OR2_X1 U592 ( .A1(G237), .A2(G902), .ZN(n498) );
  NAND2_X1 U593 ( .A1(G214), .A2(n498), .ZN(n569) );
  NAND2_X1 U594 ( .A1(G224), .A2(n736), .ZN(n492) );
  XNOR2_X1 U595 ( .A(n493), .B(n492), .ZN(n495) );
  XOR2_X1 U596 ( .A(n495), .B(n713), .Z(n496) );
  NAND2_X1 U597 ( .A1(G210), .A2(n498), .ZN(n499) );
  BUF_X2 U598 ( .A(n533), .Z(n572) );
  INV_X1 U599 ( .A(n501), .ZN(n502) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n728) );
  XOR2_X1 U601 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n505) );
  XNOR2_X1 U602 ( .A(G143), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U603 ( .A(n505), .B(n504), .ZN(n509) );
  XOR2_X1 U604 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n507) );
  XNOR2_X1 U605 ( .A(G113), .B(KEYINPUT11), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U607 ( .A(n509), .B(n508), .ZN(n514) );
  NAND2_X1 U608 ( .A1(G214), .A2(n510), .ZN(n511) );
  XNOR2_X1 U609 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U610 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U611 ( .A(n728), .B(n515), .ZN(n699) );
  NOR2_X1 U612 ( .A1(G902), .A2(n699), .ZN(n517) );
  XNOR2_X1 U613 ( .A(KEYINPUT13), .B(G475), .ZN(n516) );
  XNOR2_X1 U614 ( .A(n517), .B(n516), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n519) );
  XNOR2_X1 U616 ( .A(G116), .B(G134), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n519), .B(n518), .ZN(n522) );
  XOR2_X1 U618 ( .A(n522), .B(n521), .Z(n525) );
  NAND2_X1 U619 ( .A1(G217), .A2(n523), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n525), .B(n524), .ZN(n706) );
  INV_X1 U621 ( .A(n555), .ZN(n526) );
  NOR2_X1 U622 ( .A1(n556), .A2(n526), .ZN(n638) );
  NAND2_X1 U623 ( .A1(n526), .A2(n556), .ZN(n539) );
  INV_X1 U624 ( .A(n539), .ZN(n635) );
  NOR2_X1 U625 ( .A1(n638), .A2(n635), .ZN(n648) );
  NAND2_X1 U626 ( .A1(n648), .A2(KEYINPUT47), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n528), .B(KEYINPUT82), .ZN(n548) );
  XNOR2_X1 U628 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U630 ( .A1(n532), .A2(n538), .ZN(n560) );
  INV_X1 U631 ( .A(n569), .ZN(n653) );
  XOR2_X1 U632 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n534) );
  XNOR2_X1 U633 ( .A(KEYINPUT67), .B(n534), .ZN(n535) );
  NOR2_X1 U634 ( .A1(n560), .A2(n583), .ZN(n631) );
  XOR2_X1 U635 ( .A(n631), .B(KEYINPUT47), .Z(n537) );
  NAND2_X1 U636 ( .A1(n631), .A2(n648), .ZN(n536) );
  NAND2_X1 U637 ( .A1(n537), .A2(n536), .ZN(n546) );
  INV_X1 U638 ( .A(n576), .ZN(n605) );
  INV_X1 U639 ( .A(n605), .ZN(n664) );
  XOR2_X1 U640 ( .A(KEYINPUT6), .B(n604), .Z(n587) );
  NOR2_X1 U641 ( .A1(n539), .A2(n587), .ZN(n540) );
  NAND2_X1 U642 ( .A1(n541), .A2(n540), .ZN(n568) );
  NOR2_X1 U643 ( .A1(n568), .A2(n542), .ZN(n544) );
  XOR2_X1 U644 ( .A(KEYINPUT89), .B(KEYINPUT36), .Z(n543) );
  XNOR2_X1 U645 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U646 ( .A1(n664), .A2(n545), .ZN(n643) );
  NAND2_X1 U647 ( .A1(n546), .A2(n643), .ZN(n547) );
  NOR2_X2 U648 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U649 ( .A(n550), .B(n549), .ZN(n566) );
  XOR2_X1 U650 ( .A(n572), .B(KEYINPUT38), .Z(n649) );
  XNOR2_X1 U651 ( .A(n553), .B(n552), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n575), .A2(n635), .ZN(n554) );
  XOR2_X1 U653 ( .A(KEYINPUT41), .B(KEYINPUT112), .Z(n559) );
  NOR2_X1 U654 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U655 ( .A1(n649), .A2(n647), .ZN(n655) );
  NAND2_X1 U656 ( .A1(n655), .A2(n569), .ZN(n558) );
  XNOR2_X1 U657 ( .A(n559), .B(n558), .ZN(n674) );
  NOR2_X1 U658 ( .A1(n674), .A2(n560), .ZN(n562) );
  XNOR2_X1 U659 ( .A(KEYINPUT42), .B(KEYINPUT113), .ZN(n561) );
  XNOR2_X1 U660 ( .A(n562), .B(n561), .ZN(n745) );
  XNOR2_X1 U661 ( .A(n563), .B(KEYINPUT65), .ZN(n564) );
  XNOR2_X1 U662 ( .A(n564), .B(KEYINPUT46), .ZN(n565) );
  NOR2_X1 U663 ( .A1(n664), .A2(n568), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U665 ( .A(n571), .B(KEYINPUT43), .ZN(n573) );
  NAND2_X1 U666 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U667 ( .A(KEYINPUT108), .B(n574), .ZN(n743) );
  NAND2_X1 U668 ( .A1(n575), .A2(n638), .ZN(n645) );
  XNOR2_X1 U669 ( .A(KEYINPUT33), .B(KEYINPUT74), .ZN(n577) );
  XNOR2_X1 U670 ( .A(n578), .B(n577), .ZN(n657) );
  INV_X1 U671 ( .A(G953), .ZN(n721) );
  NOR2_X1 U672 ( .A1(G898), .A2(n721), .ZN(n716) );
  NAND2_X1 U673 ( .A1(n579), .A2(n716), .ZN(n580) );
  XOR2_X1 U674 ( .A(KEYINPUT92), .B(n580), .Z(n581) );
  NOR2_X1 U675 ( .A1(n582), .A2(n581), .ZN(n584) );
  INV_X1 U676 ( .A(n592), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n657), .A2(n594), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n586), .B(KEYINPUT88), .ZN(n600) );
  INV_X1 U679 ( .A(n587), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n604), .A2(n591), .ZN(n670) );
  NAND2_X1 U681 ( .A1(n670), .A2(n592), .ZN(n593) );
  XNOR2_X1 U682 ( .A(n593), .B(KEYINPUT31), .ZN(n639) );
  OR2_X1 U683 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U684 ( .A1(n662), .A2(n596), .ZN(n627) );
  NOR2_X1 U685 ( .A1(n639), .A2(n627), .ZN(n597) );
  NOR2_X1 U686 ( .A1(n648), .A2(n597), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n625), .A2(n598), .ZN(n599) );
  NAND2_X1 U688 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U689 ( .A(n601), .B(KEYINPUT87), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  BUF_X1 U691 ( .A(n610), .Z(n740) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT45), .ZN(n722) );
  NAND2_X1 U694 ( .A1(KEYINPUT2), .A2(n645), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT81), .B(n616), .Z(n617) );
  NAND2_X1 U696 ( .A1(G472), .A2(n708), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n624), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U698 ( .A(G101), .B(n625), .Z(G3) );
  NAND2_X1 U699 ( .A1(n627), .A2(n635), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n629) );
  NAND2_X1 U702 ( .A1(n627), .A2(n638), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U704 ( .A(G107), .B(n630), .ZN(G9) );
  XOR2_X1 U705 ( .A(G128), .B(KEYINPUT29), .Z(n633) );
  NAND2_X1 U706 ( .A1(n631), .A2(n638), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n633), .B(n632), .ZN(G30) );
  NAND2_X1 U708 ( .A1(n631), .A2(n635), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(G146), .ZN(G48) );
  NAND2_X1 U710 ( .A1(n639), .A2(n635), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT114), .ZN(n637) );
  XNOR2_X1 U712 ( .A(G113), .B(n637), .ZN(G15) );
  XOR2_X1 U713 ( .A(G116), .B(KEYINPUT115), .Z(n641) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n641), .B(n640), .ZN(G18) );
  XOR2_X1 U716 ( .A(KEYINPUT116), .B(KEYINPUT37), .Z(n642) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(G125), .B(n644), .ZN(G27) );
  XNOR2_X1 U719 ( .A(G134), .B(n645), .ZN(G36) );
  NOR2_X1 U720 ( .A1(n674), .A2(n657), .ZN(n646) );
  NOR2_X1 U721 ( .A1(G953), .A2(n646), .ZN(n689) );
  INV_X1 U722 ( .A(n647), .ZN(n651) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n677) );
  XOR2_X1 U728 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n672) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U730 ( .A(KEYINPUT49), .B(n660), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U732 ( .A(KEYINPUT118), .B(n663), .Z(n668) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U734 ( .A(KEYINPUT50), .B(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U737 ( .A(n672), .B(n671), .Z(n673) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(n675), .B(KEYINPUT120), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n678), .B(KEYINPUT52), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n687) );
  XNOR2_X1 U743 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n684) );
  NAND2_X1 U744 ( .A1(n681), .A2(n684), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT84), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n685), .A2(n362), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U748 ( .A(KEYINPUT53), .B(n690), .Z(G75) );
  NAND2_X1 U749 ( .A1(n708), .A2(G210), .ZN(n693) );
  XNOR2_X1 U750 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  NAND2_X1 U752 ( .A1(n708), .A2(G469), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n712), .A2(n698), .ZN(G54) );
  NAND2_X1 U754 ( .A1(n708), .A2(G475), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U756 ( .A(KEYINPUT60), .B(KEYINPUT68), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(G60) );
  NAND2_X1 U758 ( .A1(G478), .A2(n708), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n712), .A2(n707), .ZN(G63) );
  NAND2_X1 U761 ( .A1(G217), .A2(n708), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G66) );
  XOR2_X1 U764 ( .A(n714), .B(n713), .Z(n715) );
  XNOR2_X1 U765 ( .A(KEYINPUT123), .B(n715), .ZN(n717) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(n726) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n719) );
  NAND2_X1 U768 ( .A1(G224), .A2(G953), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(G898), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U773 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U774 ( .A(KEYINPUT122), .B(n727), .ZN(G69) );
  XNOR2_X1 U775 ( .A(n729), .B(n728), .ZN(n730) );
  XOR2_X1 U776 ( .A(n730), .B(KEYINPUT124), .Z(n735) );
  XOR2_X1 U777 ( .A(n735), .B(KEYINPUT125), .Z(n731) );
  XNOR2_X1 U778 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U779 ( .A1(G900), .A2(n732), .ZN(n733) );
  NAND2_X1 U780 ( .A1(G953), .A2(n733), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n734), .B(KEYINPUT126), .ZN(n739) );
  XNOR2_X1 U782 ( .A(n681), .B(n735), .ZN(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n739), .A2(n738), .ZN(G72) );
  XOR2_X1 U785 ( .A(G122), .B(n740), .Z(G24) );
  XOR2_X1 U786 ( .A(G119), .B(n741), .Z(G21) );
  XOR2_X1 U787 ( .A(n742), .B(G110), .Z(G12) );
  XOR2_X1 U788 ( .A(G140), .B(n743), .Z(n744) );
  XNOR2_X1 U789 ( .A(KEYINPUT117), .B(n744), .ZN(G42) );
  XNOR2_X1 U790 ( .A(G137), .B(n745), .ZN(G39) );
  XOR2_X1 U791 ( .A(G131), .B(n746), .Z(n747) );
  XNOR2_X1 U792 ( .A(KEYINPUT127), .B(n747), .ZN(G33) );
  XNOR2_X1 U793 ( .A(n748), .B(G143), .ZN(G45) );
endmodule

