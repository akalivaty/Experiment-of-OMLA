//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G155gat), .B(G162gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G155gat), .ZN(new_n208));
  INV_X1    g007(.A(G162gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT2), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G141gat), .B(G148gat), .Z(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(KEYINPUT77), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(KEYINPUT2), .C1(new_n208), .C2(new_n209), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT78), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n220), .A3(new_n206), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n213), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT73), .B(G218gat), .Z(new_n225));
  INV_X1    g024(.A(G211gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT72), .B(G197gat), .ZN(new_n228));
  INV_X1    g027(.A(G204gat), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n232), .A2(new_n234), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n223), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n222), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n235), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n239), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n223), .ZN(new_n244));
  INV_X1    g043(.A(G228gat), .ZN(new_n245));
  INV_X1    g044(.A(G233gat), .ZN(new_n246));
  OAI22_X1  g045(.A1(new_n240), .A2(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n223), .ZN(new_n248));
  INV_X1    g047(.A(new_n242), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n221), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n220), .B1(new_n217), .B2(new_n206), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n212), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n241), .B2(new_n235), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n245), .A2(new_n246), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G22gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n247), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n247), .B2(new_n257), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n205), .B(new_n259), .C1(new_n260), .C2(KEYINPUT82), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(KEYINPUT82), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n257), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(KEYINPUT81), .A3(G22gat), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n265), .A2(new_n204), .ZN(new_n266));
  INV_X1    g065(.A(new_n260), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n259), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n262), .A2(new_n263), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G113gat), .B(G120gat), .Z(new_n271));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n275), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(KEYINPUT69), .B(G127gat), .Z(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT68), .B(G134gat), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n253), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n276), .A2(new_n277), .B1(new_n284), .B2(new_n283), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n222), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G225gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT79), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n243), .A3(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(new_n292), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n288), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n296), .A2(new_n297), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n303), .A2(KEYINPUT5), .A3(new_n297), .A4(new_n296), .ZN(new_n304));
  XOR2_X1   g103(.A(G1gat), .B(G29gat), .Z(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n302), .A2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(new_n309), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT6), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n312), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(KEYINPUT65), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT24), .ZN(new_n328));
  NAND3_X1  g127(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G183gat), .B2(G190gat), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT25), .B(new_n324), .C1(new_n328), .C2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n337), .B(KEYINPUT28), .C1(new_n339), .C2(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT67), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n341), .A2(KEYINPUT26), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(KEYINPUT26), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n322), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n345), .B2(KEYINPUT66), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n338), .B(new_n346), .C1(KEYINPUT66), .C2(new_n345), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n340), .A2(new_n344), .A3(new_n325), .A4(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n336), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G226gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(new_n246), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n351), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n223), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n358));
  INV_X1    g157(.A(new_n351), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n355), .A2(new_n356), .A3(new_n242), .A4(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n360), .A2(new_n352), .A3(new_n242), .A4(new_n354), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT76), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n349), .A2(new_n351), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n359), .B1(new_n336), .B2(new_n348), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT74), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n242), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n361), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n354), .B1(new_n351), .B2(new_n349), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n367), .B1(new_n377), .B2(KEYINPUT74), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT76), .B(new_n362), .C1(new_n378), .C2(new_n242), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n361), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n270), .B1(new_n316), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT36), .ZN(new_n385));
  XOR2_X1   g184(.A(G15gat), .B(G43gat), .Z(new_n386));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n353), .A2(KEYINPUT71), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT71), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n336), .A2(new_n391), .A3(new_n348), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n286), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G227gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n394), .A2(new_n246), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n353), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n389), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT34), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(new_n396), .ZN(new_n401));
  INV_X1    g200(.A(new_n395), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI211_X1 g202(.A(KEYINPUT34), .B(new_n395), .C1(new_n393), .C2(new_n396), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n403), .A2(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(new_n399), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n413), .B2(new_n405), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n385), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n408), .B1(new_n406), .B2(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n410), .A3(new_n405), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n384), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n382), .A2(new_n381), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n380), .B1(new_n379), .B2(new_n361), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT30), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n313), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT84), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n309), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT39), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n290), .B2(new_n292), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n292), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n430), .A3(new_n292), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n436), .A2(new_n314), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT40), .B(new_n435), .C1(new_n437), .C2(new_n429), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n429), .B1(new_n436), .B2(new_n314), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n428), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT85), .B1(new_n424), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n440), .A2(new_n434), .A3(new_n439), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n314), .B1(new_n313), .B2(new_n425), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n427), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n446), .A2(new_n383), .A3(new_n447), .A4(new_n441), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n269), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n265), .A2(new_n204), .ZN(new_n451));
  INV_X1    g250(.A(new_n263), .ZN(new_n452));
  OAI22_X1  g251(.A1(new_n450), .A2(new_n451), .B1(new_n261), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n380), .C1(new_n370), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n370), .A2(new_n456), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n380), .B1(new_n370), .B2(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT86), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n454), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n380), .A2(new_n454), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n366), .A2(new_n368), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n456), .B1(new_n464), .B2(new_n242), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n355), .A2(new_n249), .A3(new_n360), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n422), .B1(new_n458), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n312), .ZN(new_n469));
  INV_X1    g268(.A(new_n427), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT84), .B1(new_n302), .B2(new_n304), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n470), .A2(new_n471), .A3(new_n314), .ZN(new_n472));
  INV_X1    g271(.A(new_n315), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n468), .B(new_n469), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n453), .B1(new_n462), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n420), .B1(new_n449), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n316), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n409), .A2(new_n414), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n453), .A2(new_n477), .A3(new_n424), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n312), .B1(new_n428), .B2(new_n315), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n481), .A2(new_n383), .A3(KEYINPUT35), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n409), .B2(new_n414), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n416), .A2(KEYINPUT87), .A3(new_n417), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n453), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n480), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  INV_X1    g289(.A(G43gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(G50gat), .ZN(new_n492));
  INV_X1    g291(.A(G50gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G43gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  AND2_X1   g296(.A1(G29gat), .A2(G36gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(KEYINPUT14), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n504));
  NAND2_X1  g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n497), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n493), .A2(G43gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n491), .A2(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n489), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT89), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT17), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n500), .A2(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT15), .B1(new_n516), .B2(new_n513), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n489), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n258), .A2(G15gat), .ZN(new_n521));
  INV_X1    g320(.A(G15gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G22gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT90), .B1(new_n527), .B2(G1gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(G8gat), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n526), .B(new_n529), .C1(KEYINPUT90), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n520), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n534), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n517), .A3(new_n519), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT18), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n534), .B(new_n532), .C1(new_n511), .C2(new_n514), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n539), .B(KEYINPUT13), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n552), .A2(new_n554), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(KEYINPUT12), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n541), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n548), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n548), .B2(new_n563), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n543), .A2(new_n547), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n568), .A2(KEYINPUT91), .B1(new_n541), .B2(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n543), .A2(new_n547), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n569), .A2(new_n571), .B1(new_n560), .B2(new_n558), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT93), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n548), .A2(new_n563), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT92), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n563), .A3(new_n564), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n568), .A2(KEYINPUT91), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n541), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n571), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n561), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n476), .A2(new_n488), .B1(new_n573), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n587), .ZN(new_n592));
  OR2_X1    g391(.A1(G57gat), .A2(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n589), .B1(new_n595), .B2(new_n585), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n601), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n535), .B1(new_n598), .B2(new_n597), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT96), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(KEYINPUT98), .A3(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  INV_X1    g423(.A(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n623), .B(new_n626), .C1(new_n591), .C2(new_n596), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n588), .A2(new_n590), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n595), .A2(new_n585), .A3(new_n589), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n618), .B1(new_n617), .B2(new_n622), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n627), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n627), .A2(new_n632), .A3(KEYINPUT101), .A4(new_n633), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n630), .A2(new_n631), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n638), .B(KEYINPUT10), .C1(new_n596), .C2(new_n591), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n612), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT103), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n612), .B1(new_n627), .B2(new_n632), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n646), .B(KEYINPUT104), .Z(new_n653));
  INV_X1    g452(.A(new_n647), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n641), .B2(new_n654), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n652), .B1(new_n651), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n607), .A2(new_n610), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n515), .B(new_n520), .C1(new_n630), .C2(new_n631), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n511), .A2(new_n514), .ZN(new_n661));
  AND2_X1   g460(.A1(G232gat), .A2(G233gat), .ZN(new_n662));
  AOI22_X1  g461(.A1(new_n661), .A2(new_n638), .B1(KEYINPUT41), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G190gat), .B(G218gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT99), .Z(new_n666));
  AND2_X1   g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n662), .A2(KEYINPUT41), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT97), .ZN(new_n671));
  XOR2_X1   g470(.A(G134gat), .B(G162gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(KEYINPUT100), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n667), .B2(new_n668), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR4_X1   g479(.A1(new_n611), .A2(new_n658), .A3(new_n659), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n584), .A2(new_n316), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n424), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n584), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT106), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(G8gat), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT107), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n687), .A2(KEYINPUT42), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n693), .B1(new_n688), .B2(new_n690), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n691), .B(new_n695), .C1(new_n696), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g496(.A1(new_n584), .A2(new_n681), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n485), .A2(new_n486), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n419), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT109), .Z(new_n706));
  AOI21_X1  g505(.A(new_n702), .B1(new_n699), .B2(new_n706), .ZN(G1326gat));
  NAND3_X1  g506(.A1(new_n699), .A2(KEYINPUT110), .A3(new_n270), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n698), .B2(new_n453), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NAND2_X1  g512(.A1(new_n384), .A2(new_n419), .ZN(new_n714));
  INV_X1    g513(.A(new_n474), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n461), .A2(new_n458), .A3(new_n457), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT38), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n270), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n443), .A2(new_n448), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n487), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n482), .B1(new_n479), .B2(KEYINPUT35), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n680), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n680), .C1(new_n720), .C2(new_n722), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n611), .A2(new_n659), .ZN(new_n728));
  INV_X1    g527(.A(new_n658), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n567), .B2(new_n572), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n577), .A2(new_n732), .A3(new_n582), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n477), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n730), .A2(new_n679), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n584), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n316), .A2(new_n502), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n740), .A2(new_n738), .A3(new_n741), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n737), .A2(new_n742), .A3(new_n743), .ZN(G1328gat));
  OAI21_X1  g543(.A(G36gat), .B1(new_n736), .B2(new_n424), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n383), .A2(new_n503), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT46), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  OR3_X1    g546(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(G1329gat));
  INV_X1    g548(.A(new_n419), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n725), .A2(new_n750), .A3(new_n726), .A4(new_n735), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n701), .A2(new_n491), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n752), .B(KEYINPUT47), .C1(new_n740), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n740), .A2(new_n753), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n727), .A2(new_n704), .A3(new_n735), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(G43gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g557(.A1(new_n725), .A2(new_n270), .A3(new_n726), .A4(new_n735), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT48), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n584), .A2(new_n493), .A3(new_n270), .A4(new_n739), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n760), .B(new_n763), .C1(new_n761), .C2(KEYINPUT48), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n728), .A2(new_n680), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n658), .A3(new_n734), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(new_n476), .B2(new_n488), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n316), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n773));
  INV_X1    g572(.A(G64gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n770), .B(new_n383), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1333gat));
  INV_X1    g576(.A(new_n770), .ZN(new_n778));
  INV_X1    g577(.A(new_n704), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(G71gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n770), .A2(new_n781), .A3(new_n701), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g583(.A1(new_n770), .A2(new_n270), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  INV_X1    g585(.A(new_n728), .ZN(new_n787));
  INV_X1    g586(.A(new_n734), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n787), .A2(new_n729), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n727), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790), .B2(new_n477), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n787), .A2(new_n788), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n680), .B(new_n792), .C1(new_n720), .C2(new_n722), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n476), .A2(new_n488), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n680), .A4(new_n792), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n316), .A2(new_n620), .A3(new_n658), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT113), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n791), .B1(new_n799), .B2(new_n801), .ZN(G1336gat));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n424), .A2(new_n729), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n621), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n424), .A2(new_n621), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n725), .A2(new_n726), .A3(new_n789), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n805), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(G92gat), .B1(new_n798), .B2(new_n806), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n814), .A2(new_n815), .A3(new_n804), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n813), .A2(new_n816), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n790), .B2(new_n779), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n700), .A2(G99gat), .A3(new_n729), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n799), .B2(new_n819), .ZN(G1338gat));
  NOR3_X1   g619(.A1(new_n453), .A2(G106gat), .A3(new_n729), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n798), .A2(new_n821), .B1(KEYINPUT116), .B2(KEYINPUT53), .ZN(new_n822));
  OR2_X1    g621(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n725), .A2(new_n270), .A3(new_n726), .A4(new_n789), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(G106gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n822), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n634), .A2(new_n635), .ZN(new_n831));
  INV_X1    g630(.A(new_n612), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n639), .A4(new_n637), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n612), .C1(new_n636), .C2(new_n640), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n646), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n830), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n642), .A2(new_n650), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n641), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n646), .A4(new_n836), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n731), .A3(new_n733), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n536), .A2(new_n538), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n540), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n545), .A2(new_n546), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n845), .A2(new_n846), .B1(new_n559), .B2(new_n555), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n567), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n658), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n680), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  INV_X1    g650(.A(new_n847), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n577), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n853), .A3(new_n680), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n848), .A2(new_n851), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n728), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n681), .A2(new_n734), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n477), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n453), .A2(new_n478), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n859), .A2(new_n424), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n788), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n857), .A2(new_n858), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n477), .A2(new_n383), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n721), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n573), .A2(new_n583), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G113gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n863), .A2(new_n869), .ZN(G1340gat));
  INV_X1    g669(.A(G120gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n866), .A2(new_n871), .A3(new_n729), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n862), .A2(new_n658), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n871), .ZN(G1341gat));
  INV_X1    g673(.A(new_n279), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n862), .A2(new_n875), .A3(new_n787), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n279), .B1(new_n866), .B2(new_n728), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  INV_X1    g677(.A(new_n281), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n879), .A3(new_n680), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT56), .Z(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n866), .B2(new_n679), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1343gat));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n865), .A2(new_n419), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n270), .A2(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(new_n849), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n573), .B2(new_n583), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n679), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n856), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n787), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n889), .B1(new_n896), .B2(new_n858), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n453), .B1(new_n857), .B2(new_n858), .ZN(new_n898));
  XNOR2_X1  g697(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n788), .B(new_n888), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G141gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n704), .A2(new_n383), .A3(new_n453), .ZN(new_n903));
  AOI21_X1  g702(.A(G141gat), .B1(new_n573), .B2(new_n583), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n859), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n887), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n887), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n867), .B(new_n888), .C1(new_n897), .C2(new_n900), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(G141gat), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT120), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(G141gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n887), .A3(new_n905), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n903), .A2(new_n859), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n901), .A2(G141gat), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n912), .B(new_n913), .C1(new_n887), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n910), .A2(new_n917), .ZN(G1344gat));
  OR2_X1    g717(.A1(new_n897), .A2(new_n900), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n658), .A4(new_n888), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n888), .A2(new_n658), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n684), .A2(new_n867), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n270), .B1(new_n923), .B2(new_n895), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n898), .A2(new_n899), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n920), .B1(new_n915), .B2(new_n658), .ZN(new_n930));
  OAI221_X1 g729(.A(new_n921), .B1(new_n928), .B2(new_n929), .C1(new_n930), .C2(G148gat), .ZN(G1345gat));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n208), .A3(new_n787), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n919), .A2(new_n888), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(new_n787), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(new_n208), .ZN(G1346gat));
  AOI21_X1  g734(.A(G162gat), .B1(new_n915), .B2(new_n680), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n679), .A2(new_n209), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n933), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n424), .A2(new_n316), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n857), .B2(new_n858), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n942), .A2(new_n860), .ZN(new_n943));
  AOI21_X1  g742(.A(G169gat), .B1(new_n943), .B2(new_n788), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n942), .A2(new_n487), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n317), .B1(new_n573), .B2(new_n583), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1348gat));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n318), .A3(new_n658), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n942), .A2(new_n487), .A3(new_n729), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n318), .B2(new_n949), .ZN(G1349gat));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n728), .A2(new_n339), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n941), .A2(new_n861), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G183gat), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n864), .A2(new_n721), .A3(new_n787), .A4(new_n939), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(KEYINPUT121), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n941), .A2(new_n957), .A3(new_n721), .A4(new_n787), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n953), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT60), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g762(.A(KEYINPUT122), .B(new_n953), .C1(new_n956), .C2(new_n958), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n955), .A2(KEYINPUT121), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(G183gat), .A3(new_n958), .ZN(new_n967));
  INV_X1    g766(.A(new_n953), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n959), .A2(new_n962), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(new_n971), .A3(new_n951), .A4(KEYINPUT60), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n965), .A2(new_n972), .ZN(G1350gat));
  INV_X1    g772(.A(G190gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n943), .A2(new_n974), .A3(new_n680), .ZN(new_n975));
  INV_X1    g774(.A(new_n945), .ZN(new_n976));
  OAI21_X1  g775(.A(G190gat), .B1(new_n976), .B2(new_n679), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n977), .A2(KEYINPUT61), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G1351gat));
  NAND2_X1  g779(.A1(new_n779), .A2(new_n939), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n981), .B1(new_n926), .B2(new_n927), .ZN(new_n982));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n983), .B1(new_n573), .B2(new_n583), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n704), .A2(new_n453), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n985), .A2(new_n788), .A3(new_n941), .ZN(new_n986));
  AOI22_X1  g785(.A1(new_n982), .A2(new_n984), .B1(new_n983), .B2(new_n986), .ZN(G1352gat));
  NAND4_X1  g786(.A1(new_n985), .A2(new_n229), .A3(new_n658), .A4(new_n941), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n229), .B1(new_n982), .B2(new_n658), .ZN(new_n990));
  OR3_X1    g789(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT124), .ZN(new_n991));
  OAI21_X1  g790(.A(KEYINPUT124), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n985), .A2(new_n226), .A3(new_n787), .A4(new_n941), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n982), .A2(new_n787), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  NAND3_X1  g797(.A1(new_n985), .A2(new_n680), .A3(new_n941), .ZN(new_n999));
  INV_X1    g798(.A(G218gat), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g800(.A1(new_n1001), .A2(KEYINPUT125), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(KEYINPUT125), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n982), .A2(KEYINPUT126), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n679), .A2(new_n225), .ZN(new_n1005));
  XNOR2_X1  g804(.A(new_n1005), .B(KEYINPUT127), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1006), .B1(new_n982), .B2(KEYINPUT126), .ZN(new_n1007));
  AOI22_X1  g806(.A1(new_n1002), .A2(new_n1003), .B1(new_n1004), .B2(new_n1007), .ZN(G1355gat));
endmodule


