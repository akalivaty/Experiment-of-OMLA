//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999;
  XOR2_X1   g000(.A(G169gat), .B(G197gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G113gat), .B(G141gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT94), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n204), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT12), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n209), .A2(KEYINPUT16), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n211), .A2(G8gat), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n209), .A2(new_n210), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(KEYINPUT16), .A3(new_n210), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n230), .A2(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT15), .ZN(new_n232));
  XOR2_X1   g031(.A(G43gat), .B(G50gat), .Z(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT17), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(KEYINPUT15), .A3(new_n233), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n219), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT95), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n219), .B(KEYINPUT95), .C1(new_n238), .C2(new_n239), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT96), .B1(new_n213), .B2(new_n217), .ZN(new_n245));
  OAI21_X1  g044(.A(G8gat), .B1(new_n211), .B2(new_n212), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT96), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n215), .A2(new_n214), .A3(new_n216), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n245), .A2(new_n249), .B1(new_n237), .B2(new_n235), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n242), .A2(new_n243), .A3(new_n244), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n208), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n237), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT17), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n218), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n250), .B1(new_n260), .B2(KEYINPUT95), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n242), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n249), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(new_n257), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n243), .B(KEYINPUT13), .Z(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n254), .A2(new_n262), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n253), .B1(new_n264), .B2(new_n265), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT97), .B1(new_n252), .B2(new_n253), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n269), .B(new_n262), .C1(new_n270), .C2(new_n208), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n274));
  XNOR2_X1  g073(.A(G127gat), .B(G134gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G113gat), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  NAND2_X1  g080(.A1(G113gat), .A2(G120gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n277), .A2(KEYINPUT70), .A3(new_n283), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n281), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n280), .A2(new_n282), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n293), .A2(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT83), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n288), .A2(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT83), .ZN(new_n301));
  XOR2_X1   g100(.A(G141gat), .B(G148gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G155gat), .B(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(KEYINPUT2), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n309), .A2(new_n308), .A3(KEYINPUT2), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n302), .B(new_n305), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n299), .A2(new_n301), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n274), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n313), .A2(KEYINPUT84), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n312), .A3(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n300), .A2(KEYINPUT4), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n326), .A3(new_n318), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT82), .B1(new_n313), .B2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n307), .A2(new_n330), .A3(new_n312), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n313), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n299), .A2(new_n332), .A3(new_n301), .A4(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT85), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  AND4_X1   g134(.A1(new_n299), .A2(new_n332), .A3(new_n301), .A4(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n336), .A2(new_n327), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n320), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n325), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n321), .B1(new_n340), .B2(new_n297), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n334), .B(new_n341), .C1(new_n321), .C2(new_n316), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n318), .A2(new_n274), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT0), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n339), .A2(new_n350), .A3(new_n345), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n328), .A2(KEYINPUT85), .A3(new_n334), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n337), .B1(new_n336), .B2(new_n327), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n344), .B1(new_n358), .B2(new_n320), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n350), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n363));
  INV_X1    g162(.A(G169gat), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT26), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n367), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n365), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n369), .A2(new_n373), .B1(G183gat), .B2(G190gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(KEYINPUT28), .A3(new_n376), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n374), .A2(KEYINPUT68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(KEYINPUT68), .B2(new_n374), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n370), .A2(KEYINPUT23), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n372), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n366), .A2(KEYINPUT23), .A3(new_n368), .ZN(new_n386));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n386), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT66), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT66), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n385), .A2(new_n386), .A3(new_n392), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n390), .B(new_n391), .C1(new_n398), .C2(KEYINPUT64), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(KEYINPUT64), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n372), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT23), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n372), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n383), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n382), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n362), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G211gat), .A2(G218gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT76), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT76), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G204gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G197gat), .ZN(new_n418));
  INV_X1    g217(.A(G197gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(G204gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n418), .B(new_n420), .C1(new_n421), .C2(KEYINPUT22), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT77), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT77), .B(new_n422), .C1(new_n414), .C2(new_n415), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n408), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n408), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n362), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n397), .A2(new_n404), .A3(KEYINPUT67), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n382), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT67), .B1(new_n397), .B2(new_n404), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n407), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n431), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n433), .A2(new_n434), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(KEYINPUT29), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n362), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n437), .B(new_n429), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(KEYINPUT80), .A3(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n445), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n441), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(KEYINPUT30), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n361), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457));
  NAND2_X1  g256(.A1(G228gat), .A2(G233gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n439), .B1(new_n313), .B2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g258(.A(new_n428), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n426), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n411), .A2(new_n412), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n464), .A2(new_n413), .A3(new_n422), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n422), .B1(new_n464), .B2(new_n413), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n439), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n330), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n340), .A2(new_n468), .A3(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n461), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT86), .B1(new_n340), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT87), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n429), .A2(new_n474), .A3(new_n459), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n424), .A2(new_n425), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n330), .B1(new_n476), .B2(KEYINPUT29), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n458), .B1(new_n477), .B2(new_n313), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G22gat), .ZN(new_n480));
  XOR2_X1   g279(.A(G78gat), .B(G106gat), .Z(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G50gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n472), .A2(new_n479), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n480), .B1(new_n472), .B2(new_n479), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n479), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(G22gat), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n485), .B2(new_n486), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n457), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n487), .A2(new_n488), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n485), .A3(new_n486), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT89), .A4(new_n484), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n300), .B1(new_n433), .B2(new_n434), .ZN(new_n499));
  INV_X1    g298(.A(G227gat), .ZN(new_n500));
  INV_X1    g299(.A(G233gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n405), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n504), .A2(new_n297), .A3(new_n432), .A4(new_n382), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n505), .A3(KEYINPUT72), .A4(new_n502), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT74), .ZN(new_n512));
  XOR2_X1   g311(.A(G71gat), .B(G99gat), .Z(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(KEYINPUT73), .B(KEYINPUT33), .Z(new_n516));
  OAI21_X1  g315(.A(KEYINPUT32), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n498), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT75), .B(new_n517), .C1(new_n508), .C2(new_n509), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n508), .B2(new_n509), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n519), .A2(new_n520), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n499), .A2(new_n505), .ZN(new_n524));
  INV_X1    g323(.A(new_n502), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n526), .A2(KEYINPUT34), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(KEYINPUT34), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  OAI221_X1 g330(.A(new_n529), .B1(new_n515), .B2(new_n522), .C1(new_n519), .C2(new_n520), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR3_X1   g332(.A1(new_n456), .A2(new_n497), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n454), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT90), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT6), .B1(new_n359), .B2(new_n350), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n350), .B(KEYINPUT91), .Z(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n359), .B2(KEYINPUT92), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n339), .A2(KEYINPUT92), .A3(new_n345), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n352), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT35), .B1(new_n493), .B2(new_n496), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n534), .A2(new_n535), .B1(new_n533), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n442), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT37), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n451), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n551), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT38), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n438), .A2(new_n440), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n431), .B2(new_n406), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n556), .B2(new_n430), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n407), .A2(new_n429), .A3(new_n435), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT38), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n559), .A2(new_n552), .B1(new_n550), .B2(new_n451), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n545), .A2(new_n554), .A3(new_n560), .A4(new_n352), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n493), .A2(new_n496), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n543), .A2(new_n544), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT39), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n342), .A2(new_n564), .A3(new_n319), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n342), .A2(new_n319), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT39), .B1(new_n317), .B2(new_n319), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n541), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT40), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n561), .B(new_n562), .C1(new_n570), .C2(new_n539), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n531), .A2(new_n572), .A3(new_n532), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n531), .B2(new_n532), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n456), .A2(new_n497), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n273), .B1(new_n549), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(KEYINPUT102), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT8), .ZN(new_n587));
  INV_X1    g386(.A(G85gat), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n583), .A2(new_n585), .A3(new_n587), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(new_n592), .A3(new_n583), .A4(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n238), .B2(new_n239), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT103), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n600), .B(new_n597), .C1(new_n238), .C2(new_n239), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n597), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n257), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G232gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(new_n501), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n580), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n609), .A3(new_n580), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT104), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n579), .B(new_n608), .C1(new_n599), .C2(new_n601), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n614), .B(new_n621), .C1(new_n610), .C2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(G71gat), .A2(G78gat), .ZN(new_n628));
  OR2_X1    g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G57gat), .A2(G64gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(G57gat), .A2(G64gat), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(G57gat), .ZN(new_n637));
  INV_X1    g436(.A(G64gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n636), .B1(new_n639), .B2(new_n632), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n631), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n639), .A2(KEYINPUT9), .A3(new_n632), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n629), .A2(KEYINPUT98), .ZN(new_n643));
  OR3_X1    g442(.A1(KEYINPUT98), .A2(G71gat), .A3(G78gat), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n628), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n245), .B(new_n249), .C1(new_n627), .C2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n627), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n627), .A3(new_n652), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n656), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n650), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n650), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n649), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n649), .B1(new_n660), .B2(new_n663), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n626), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n649), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n660), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n664), .A3(new_n625), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n623), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n646), .A2(new_n597), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n641), .A2(new_n594), .A3(new_n645), .A4(new_n596), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n645), .A4(new_n641), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n680), .B2(new_n682), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n679), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n686), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n683), .B2(new_n684), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n688), .A3(new_n678), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n675), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n687), .A2(new_n689), .A3(new_n679), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n678), .B1(new_n692), .B2(new_n688), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n578), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n361), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n210), .ZN(G1324gat));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(new_n539), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT42), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n704), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(G8gat), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n707), .B2(new_n711), .ZN(G1325gat));
  OAI21_X1  g511(.A(G15gat), .B1(new_n701), .B2(new_n575), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n533), .A2(G15gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n701), .B2(new_n714), .ZN(G1326gat));
  NAND3_X1  g514(.A1(new_n704), .A2(KEYINPUT107), .A3(new_n497), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n701), .B2(new_n562), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  NOR3_X1   g520(.A1(new_n623), .A2(new_n673), .A3(new_n698), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n578), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n361), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n228), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n549), .A2(new_n577), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n623), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n667), .A2(new_n732), .A3(new_n671), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n667), .B2(new_n671), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n273), .A3(new_n698), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n346), .A2(new_n351), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n540), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n454), .B1(new_n738), .B2(new_n352), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n739), .B2(new_n562), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n456), .A2(new_n497), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n575), .A3(new_n571), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n623), .B1(new_n744), .B2(new_n549), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n731), .B(new_n736), .C1(new_n745), .C2(KEYINPUT44), .ZN(new_n746));
  OAI21_X1  g545(.A(G29gat), .B1(new_n746), .B2(new_n361), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n747), .ZN(G1328gat));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n539), .A2(G36gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n578), .A2(new_n749), .A3(new_n722), .A4(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT110), .Z(new_n752));
  OAI21_X1  g551(.A(G36gat), .B1(new_n746), .B2(new_n539), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n723), .A2(G36gat), .A3(new_n539), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n752), .B(new_n753), .C1(new_n749), .C2(new_n754), .ZN(G1329gat));
  NOR2_X1   g554(.A1(new_n723), .A2(new_n533), .ZN(new_n756));
  INV_X1    g555(.A(new_n575), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  OAI22_X1  g557(.A1(G43gat), .A2(new_n756), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n549), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n620), .A2(new_n622), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n764), .A2(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(KEYINPUT111), .A3(new_n497), .A4(new_n736), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n746), .B2(new_n562), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n562), .A2(G50gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n724), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT48), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n729), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n497), .A3(new_n731), .A4(new_n736), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n774), .A2(G50gat), .B1(new_n724), .B2(new_n770), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n769), .A2(new_n772), .B1(KEYINPUT48), .B2(new_n775), .ZN(G1331gat));
  INV_X1    g575(.A(new_n698), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n674), .A2(new_n272), .A3(new_n777), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n762), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n725), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g580(.A1(new_n779), .A2(new_n705), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT49), .B(G64gat), .Z(new_n783));
  AND2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT112), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n783), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n788), .B(new_n789), .C1(new_n785), .C2(new_n782), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1333gat));
  NAND3_X1  g590(.A1(new_n779), .A2(G71gat), .A3(new_n757), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n533), .B(KEYINPUT113), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n795), .B2(G71gat), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n497), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g598(.A1(new_n673), .A2(new_n272), .A3(new_n777), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n731), .B(new_n800), .C1(new_n745), .C2(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801), .B2(new_n361), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n673), .A2(new_n272), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n762), .A2(new_n763), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n725), .A2(new_n588), .A3(new_n698), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n802), .B1(new_n809), .B2(new_n810), .ZN(G1336gat));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n765), .A2(new_n812), .A3(new_n705), .A4(new_n800), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT114), .B1(new_n801), .B2(new_n539), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n589), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n539), .A2(G92gat), .A3(new_n777), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n773), .A2(new_n705), .A3(new_n731), .A4(new_n800), .ZN(new_n820));
  AOI22_X1  g619(.A1(G92gat), .A2(new_n820), .B1(new_n808), .B2(new_n816), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n815), .A2(new_n819), .B1(new_n821), .B2(new_n818), .ZN(G1337gat));
  OAI21_X1  g621(.A(KEYINPUT115), .B1(new_n801), .B2(new_n575), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G99gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n575), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n533), .A2(G99gat), .A3(new_n777), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT116), .Z(new_n827));
  OAI22_X1  g626(.A1(new_n824), .A2(new_n825), .B1(new_n809), .B2(new_n827), .ZN(G1338gat));
  NOR3_X1   g627(.A1(new_n562), .A2(G106gat), .A3(new_n777), .ZN(new_n829));
  INV_X1    g628(.A(new_n807), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT51), .B1(new_n745), .B2(new_n803), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G106gat), .B1(new_n801), .B2(new_n562), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1339gat));
  NAND3_X1  g637(.A1(new_n683), .A2(new_n684), .A3(new_n691), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n687), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n679), .B1(new_n692), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n695), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n683), .A2(new_n684), .A3(new_n691), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n692), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n685), .A2(new_n841), .A3(new_n686), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n678), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT117), .B(new_n845), .C1(new_n847), .C2(new_n849), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n844), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n271), .B2(new_n268), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n254), .A2(new_n208), .A3(new_n262), .A4(new_n266), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n243), .B1(new_n261), .B2(new_n242), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n264), .A2(new_n265), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n207), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n856), .A2(new_n698), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n623), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n844), .A2(new_n852), .A3(new_n853), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n856), .A2(new_n859), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n620), .A2(new_n862), .A3(new_n863), .A4(new_n622), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n735), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n273), .A2(new_n623), .A3(new_n673), .A4(new_n777), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT118), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n860), .B1(new_n272), .B2(new_n862), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n869), .B2(new_n763), .ZN(new_n870));
  INV_X1    g669(.A(new_n735), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n866), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n705), .A2(new_n361), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n868), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n497), .A2(new_n533), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n273), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(new_n278), .ZN(G1340gat));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n777), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n279), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n878), .B2(new_n871), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n672), .A2(G127gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n878), .B2(new_n884), .ZN(G1342gat));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n877), .A3(new_n763), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G134gat), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(G134gat), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n889), .A2(KEYINPUT119), .A3(new_n888), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n889), .B2(new_n888), .ZN(new_n891));
  OAI221_X1 g690(.A(new_n887), .B1(new_n888), .B2(new_n889), .C1(new_n890), .C2(new_n891), .ZN(G1343gat));
  NAND3_X1  g691(.A1(new_n868), .A2(new_n874), .A3(new_n497), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n844), .A2(new_n850), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n268), .B2(new_n271), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n623), .B1(new_n897), .B2(new_n860), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT120), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n623), .B(new_n900), .C1(new_n897), .C2(new_n860), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(new_n864), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n866), .B1(new_n902), .B2(new_n673), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n562), .A2(new_n894), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n875), .A2(new_n575), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n272), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n573), .A2(new_n574), .A3(new_n562), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n868), .A2(new_n874), .A3(new_n912), .A4(new_n875), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n273), .A2(G141gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n910), .B(new_n911), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n876), .A2(KEYINPUT121), .A3(new_n912), .A4(new_n914), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n913), .B2(new_n915), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n917), .B(new_n911), .C1(new_n910), .C2(new_n921), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n893), .A2(new_n894), .B1(new_n903), .B2(new_n904), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n273), .A3(new_n907), .ZN(new_n924));
  INV_X1    g723(.A(G141gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT122), .B1(new_n926), .B2(KEYINPUT58), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n916), .B1(new_n922), .B2(new_n927), .ZN(G1344gat));
  INV_X1    g727(.A(new_n913), .ZN(new_n929));
  INV_X1    g728(.A(G148gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(new_n698), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n923), .A2(new_n907), .ZN(new_n932));
  AOI211_X1 g731(.A(KEYINPUT59), .B(new_n930), .C1(new_n932), .C2(new_n698), .ZN(new_n933));
  XOR2_X1   g732(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n934));
  AND2_X1   g733(.A1(new_n700), .A2(new_n273), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n673), .B1(new_n898), .B2(new_n864), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n894), .B(new_n497), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n698), .A4(new_n908), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n934), .B1(new_n939), .B2(G148gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n931), .B1(new_n933), .B2(new_n940), .ZN(G1345gat));
  NOR2_X1   g740(.A1(new_n913), .A2(new_n672), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT124), .ZN(new_n943));
  AOI21_X1  g742(.A(G155gat), .B1(new_n942), .B2(KEYINPUT124), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n735), .A2(G155gat), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n943), .A2(new_n944), .B1(new_n932), .B2(new_n945), .ZN(G1346gat));
  INV_X1    g745(.A(G162gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n947), .A3(new_n763), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n923), .A2(new_n623), .A3(new_n907), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n947), .ZN(G1347gat));
  AND2_X1   g749(.A1(new_n868), .A2(new_n874), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n539), .A2(new_n725), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n951), .A2(new_n877), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n272), .A2(new_n364), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n951), .A2(new_n562), .A3(new_n794), .A4(new_n952), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n273), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n953), .B2(new_n955), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT126), .ZN(G1348gat));
  OAI21_X1  g760(.A(G176gat), .B1(new_n957), .B2(new_n777), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n698), .A2(new_n365), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n953), .B2(new_n963), .ZN(G1349gat));
  INV_X1    g763(.A(new_n953), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n375), .A3(new_n673), .ZN(new_n966));
  OAI21_X1  g765(.A(G183gat), .B1(new_n957), .B2(new_n871), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n376), .A3(new_n763), .ZN(new_n970));
  OAI21_X1  g769(.A(G190gat), .B1(new_n957), .B2(new_n623), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n973), .B(G190gat), .C1(new_n957), .C2(new_n623), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n975), .B2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n970), .B1(new_n976), .B2(new_n978), .ZN(G1351gat));
  NAND3_X1  g778(.A1(new_n951), .A2(new_n912), .A3(new_n952), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n272), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n937), .A2(new_n938), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n575), .A2(new_n952), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n273), .A2(new_n419), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n982), .B1(new_n985), .B2(new_n986), .ZN(G1352gat));
  NOR3_X1   g786(.A1(new_n980), .A2(G204gat), .A3(new_n777), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n983), .A2(new_n777), .A3(new_n984), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n417), .B2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n981), .A2(new_n409), .A3(new_n673), .ZN(new_n992));
  INV_X1    g791(.A(new_n984), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n937), .A2(new_n938), .A3(new_n673), .A4(new_n993), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n994), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n994), .B2(G211gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G1354gat));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n410), .A3(new_n763), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n983), .A2(new_n623), .A3(new_n984), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n410), .ZN(G1355gat));
endmodule


