//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G125), .B(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(KEYINPUT16), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(G146), .A3(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n200), .A2(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n203), .C1(new_n204), .C2(KEYINPUT23), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  XNOR2_X1  g020(.A(G119), .B(G128), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n199), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n191), .A2(KEYINPUT76), .A3(new_n194), .A4(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n190), .A2(new_n196), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT75), .B(G110), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n205), .A2(new_n214), .B1(new_n206), .B2(new_n207), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G953), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(G221), .A3(G234), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT77), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G137), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n209), .B2(new_n216), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT25), .B1(new_n226), .B2(new_n188), .ZN(new_n227));
  OAI211_X1 g041(.A(KEYINPUT25), .B(new_n188), .C1(new_n224), .C2(new_n225), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n189), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n226), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n189), .A2(G902), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n196), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n236), .A2(G146), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n196), .A2(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n239), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT0), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(KEYINPUT0), .B2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n247), .A2(new_n249), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n235), .A2(new_n237), .B1(KEYINPUT0), .B2(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT65), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n241), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G134), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G137), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n258), .B1(KEYINPUT11), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT11), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n259), .B2(G137), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(G131), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n245), .B1(new_n244), .B2(new_n250), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT65), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n240), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n256), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n242), .A2(new_n243), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n202), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n260), .B2(new_n258), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n276), .B(new_n277), .C1(G131), .C2(new_n264), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(KEYINPUT2), .A2(G113), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT66), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(KEYINPUT2), .B2(G113), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n281), .A2(new_n283), .B1(KEYINPUT2), .B2(G113), .ZN(new_n284));
  XNOR2_X1  g098(.A(G116), .B(G119), .ZN(new_n285));
  AOI211_X1 g099(.A(KEYINPUT67), .B(KEYINPUT68), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n283), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT2), .A2(G113), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n285), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n286), .A2(new_n292), .B1(new_n284), .B2(new_n285), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n291), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n284), .A2(new_n285), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(new_n291), .A3(new_n287), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n279), .A2(KEYINPUT72), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n271), .A2(new_n299), .A3(new_n278), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n271), .A2(new_n299), .A3(KEYINPUT28), .A4(new_n278), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n279), .B2(new_n299), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n300), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G210), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n310), .B(KEYINPUT27), .Z(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G101), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n311), .B(new_n312), .Z(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(KEYINPUT29), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n303), .A2(new_n304), .ZN(new_n317));
  INV_X1    g131(.A(new_n299), .ZN(new_n318));
  INV_X1    g132(.A(G131), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n264), .B(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n278), .B1(new_n320), .B2(new_n255), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n317), .A2(KEYINPUT71), .A3(new_n313), .A4(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT71), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n303), .A2(new_n322), .A3(new_n304), .ZN(new_n325));
  INV_X1    g139(.A(new_n313), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n271), .A2(KEYINPUT30), .A3(new_n278), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n318), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n301), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n332), .B2(new_n326), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n323), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n308), .A2(new_n335), .A3(new_n314), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n316), .A2(new_n334), .A3(new_n188), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G472), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(KEYINPUT74), .A3(G472), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n331), .A2(new_n313), .A3(new_n301), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT31), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n325), .A2(new_n326), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n331), .A2(new_n346), .A3(new_n313), .A4(new_n301), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT70), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(KEYINPUT70), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n234), .B1(new_n342), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G469), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n188), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n362), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G107), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G101), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n368), .A2(G101), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n363), .A2(new_n366), .A3(new_n372), .A4(new_n367), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT79), .B(new_n370), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(G101), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT4), .A4(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n256), .A2(new_n379), .A3(new_n270), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT80), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n256), .A2(new_n379), .A3(KEYINPUT80), .A4(new_n270), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND4_X1   g198(.A1(new_n273), .A2(new_n235), .A3(new_n237), .A4(G128), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT81), .B1(new_n242), .B2(new_n273), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n235), .A2(new_n387), .A3(KEYINPUT1), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G128), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n385), .B1(new_n389), .B2(new_n238), .ZN(new_n390));
  INV_X1    g204(.A(new_n367), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n362), .A2(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n373), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n394), .A2(KEYINPUT82), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(KEYINPUT82), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n276), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n395), .B1(KEYINPUT10), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n384), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n265), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n218), .A2(G227), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT78), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n266), .A2(new_n267), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n269), .B1(new_n407), .B2(new_n241), .ZN(new_n408));
  AOI211_X1 g222(.A(KEYINPUT69), .B(new_n240), .C1(new_n266), .C2(new_n267), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT80), .B1(new_n410), .B2(new_n379), .ZN(new_n411));
  AND4_X1   g225(.A1(KEYINPUT80), .A2(new_n256), .A3(new_n379), .A4(new_n270), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n320), .B(new_n400), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n406), .A3(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n390), .A2(new_n394), .ZN(new_n415));
  INV_X1    g229(.A(new_n394), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n276), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n265), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n418), .B(KEYINPUT12), .Z(new_n419));
  AOI21_X1  g233(.A(new_n406), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT83), .B(new_n361), .C1(new_n422), .C2(new_n359), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n320), .B1(new_n384), .B2(new_n400), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n265), .B(new_n399), .C1(new_n382), .C2(new_n383), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n420), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n424), .B(G469), .C1(new_n428), .C2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n406), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n425), .B2(new_n426), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n413), .A2(KEYINPUT84), .A3(new_n406), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n419), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT84), .B1(new_n413), .B2(new_n406), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n359), .A3(new_n188), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(G952), .A3(new_n218), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(G898), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G214), .B1(G237), .B2(G902), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n293), .A2(new_n298), .A3(new_n379), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n200), .A2(G116), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n446), .B(G113), .C1(KEYINPUT5), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n290), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n397), .A3(new_n396), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G122), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n451), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G125), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n274), .B(new_n458), .C1(new_n272), .C2(new_n275), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n268), .A2(new_n458), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT85), .B1(new_n268), .B2(new_n458), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G224), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G953), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n467), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n463), .A2(new_n469), .A3(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n452), .A2(new_n472), .A3(new_n454), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n457), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n459), .B1(new_n268), .B2(new_n458), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n469), .A2(KEYINPUT7), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n450), .A2(new_n394), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n453), .B(KEYINPUT8), .Z(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n449), .B2(new_n416), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n475), .A2(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n456), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n476), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n463), .A2(KEYINPUT86), .A3(new_n464), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n255), .A2(new_n462), .A3(G125), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(new_n464), .A3(new_n459), .A4(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n474), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n474), .B2(new_n489), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n443), .B(new_n444), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n236), .A2(G128), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n202), .A2(G143), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G134), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n259), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT92), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n504));
  INV_X1    g318(.A(G122), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(G116), .ZN(new_n506));
  INV_X1    g320(.A(G116), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(KEYINPUT89), .A3(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT14), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(G116), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n509), .A2(KEYINPUT14), .ZN(new_n513));
  OAI21_X1  g327(.A(G107), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n365), .A3(new_n511), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n503), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n494), .B2(new_n517), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT90), .B(KEYINPUT13), .C1(new_n236), .C2(G128), .ZN(new_n520));
  OAI221_X1 g334(.A(new_n495), .B1(new_n517), .B2(new_n494), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G134), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n511), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G107), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n515), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n498), .B(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT9), .B(G234), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n528), .A2(new_n187), .A3(G953), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n516), .B2(new_n527), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n188), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G478), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n533), .B(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G475), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(G143), .B1(new_n309), .B2(G214), .ZN(new_n541));
  OAI21_X1  g355(.A(G131), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n309), .A2(G214), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n236), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n319), .A3(new_n539), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT17), .B(G131), .C1(new_n540), .C2(new_n541), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n197), .A3(new_n198), .A4(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT88), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(G104), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(G104), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n556), .A2(KEYINPUT88), .A3(new_n552), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n539), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT18), .A2(G131), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n458), .A2(G140), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n193), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G146), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n559), .A2(new_n561), .B1(new_n565), .B2(new_n213), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n549), .A2(new_n558), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n549), .A2(new_n567), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n556), .A2(new_n552), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n538), .B1(new_n571), .B2(new_n188), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n542), .A2(new_n545), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n190), .A2(KEYINPUT19), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n190), .A2(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n196), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n211), .A2(new_n573), .A3(new_n576), .A4(new_n212), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n567), .ZN(new_n578));
  INV_X1    g392(.A(new_n570), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n568), .ZN(new_n581));
  NOR2_X1   g395(.A1(G475), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT20), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT20), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n585), .A3(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n572), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n537), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n493), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G221), .B1(new_n528), .B2(G902), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n437), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n358), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT93), .B(G101), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G3));
  AND2_X1   g408(.A1(new_n437), .A2(new_n590), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n348), .A2(new_n188), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n350), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n234), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n493), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n534), .A2(new_n188), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n516), .A2(new_n527), .ZN(new_n603));
  INV_X1    g417(.A(new_n529), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(G902), .B1(new_n605), .B2(new_n530), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n606), .B2(new_n534), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n531), .B2(new_n532), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n605), .A2(new_n609), .A3(new_n530), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n610), .A3(G478), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n587), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n600), .A2(new_n601), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  AOI21_X1  g430(.A(new_n585), .B1(new_n581), .B2(new_n582), .ZN(new_n617));
  INV_X1    g431(.A(new_n582), .ZN(new_n618));
  AOI211_X1 g432(.A(KEYINPUT20), .B(new_n618), .C1(new_n580), .C2(new_n568), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n572), .B1(new_n621), .B2(KEYINPUT94), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(new_n537), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n600), .A2(new_n601), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n217), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n232), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n230), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n598), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n635), .A2(new_n590), .A3(new_n437), .A4(new_n589), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT37), .B(G110), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  AND3_X1   g452(.A1(new_n337), .A2(KEYINPUT74), .A3(G472), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT74), .B1(new_n337), .B2(G472), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n357), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n444), .B(new_n633), .C1(new_n491), .C2(new_n492), .ZN(new_n642));
  INV_X1    g456(.A(new_n439), .ZN(new_n643));
  INV_X1    g457(.A(new_n440), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(G900), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n622), .A2(new_n536), .A3(new_n624), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n437), .A2(new_n647), .A3(new_n590), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n645), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n595), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n492), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n474), .A2(new_n489), .A3(new_n490), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n568), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n570), .B1(new_n549), .B2(new_n567), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n188), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G475), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n617), .B2(new_n619), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n536), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n634), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n444), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n332), .A2(new_n313), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n307), .B(new_n301), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n188), .B(new_n671), .C1(new_n672), .C2(new_n313), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G472), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n357), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n670), .B1(new_n357), .B2(new_n674), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n659), .B(new_n669), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n654), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n236), .ZN(G45));
  INV_X1    g496(.A(new_n612), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n664), .A4(new_n645), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n664), .A2(new_n611), .A3(new_n607), .A4(new_n645), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n642), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n689), .A2(new_n437), .A3(new_n590), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n641), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NAND2_X1  g506(.A1(new_n435), .A2(new_n188), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n590), .A3(new_n436), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n695), .A2(new_n493), .A3(new_n587), .A4(new_n612), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n358), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NOR4_X1   g513(.A1(new_n695), .A2(new_n493), .A3(new_n537), .A4(new_n625), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n358), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  NOR4_X1   g516(.A1(new_n695), .A2(new_n442), .A3(new_n588), .A4(new_n642), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n641), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND2_X1  g519(.A1(new_n694), .A2(new_n436), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n344), .B(new_n347), .C1(new_n308), .C2(new_n313), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n349), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n597), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n234), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n493), .A2(new_n665), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n711), .A3(new_n590), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  AOI21_X1  g528(.A(new_n668), .B1(new_n655), .B2(new_n656), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n694), .A2(new_n590), .A3(new_n436), .A4(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n685), .A2(new_n687), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n597), .A3(new_n633), .A4(new_n709), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT99), .B(G125), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G27));
  INV_X1    g535(.A(KEYINPUT84), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n426), .B2(new_n430), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n419), .A3(new_n432), .ZN(new_n724));
  AOI21_X1  g538(.A(G902), .B1(new_n724), .B2(new_n431), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n360), .B1(new_n725), .B2(new_n359), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT100), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n414), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(G469), .B(new_n728), .C1(new_n428), .C2(new_n727), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n422), .A2(KEYINPUT100), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT101), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n732), .A3(G469), .A4(new_n728), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n726), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n590), .A2(new_n444), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n657), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n734), .A2(KEYINPUT102), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT102), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n717), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n354), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT32), .B1(new_n348), .B2(new_n349), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n234), .B1(new_n342), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT42), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n688), .A2(KEYINPUT42), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n358), .B(new_n747), .C1(new_n738), .C2(new_n737), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n319), .ZN(G33));
  INV_X1    g564(.A(new_n646), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n358), .B(new_n751), .C1(new_n738), .C2(new_n737), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NOR2_X1   g567(.A1(new_n657), .A2(new_n668), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n634), .B1(new_n597), .B2(new_n350), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n612), .A2(new_n664), .A3(KEYINPUT43), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n612), .B1(new_n758), .B2(new_n664), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n664), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n757), .B1(new_n760), .B2(KEYINPUT43), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n755), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT44), .B(new_n756), .C1(new_n762), .C2(new_n763), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n359), .B1(new_n422), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n728), .B1(new_n428), .B2(new_n727), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT46), .A3(new_n361), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT104), .A3(new_n436), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n774), .A2(new_n361), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n776), .B1(KEYINPUT46), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT104), .B1(new_n775), .B2(new_n436), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n590), .B(new_n651), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n769), .A2(new_n770), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n257), .ZN(G39));
  AOI22_X1  g596(.A1(new_n340), .A2(new_n341), .B1(new_n356), .B2(new_n355), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n234), .A3(new_n717), .A4(new_n754), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n590), .B1(new_n778), .B2(new_n779), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n192), .ZN(G42));
  NOR2_X1   g604(.A1(G952), .A2(G953), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT119), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n787), .B(new_n788), .C1(new_n590), .C2(new_n706), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n711), .A2(new_n439), .A3(new_n761), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n754), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n695), .A2(new_n444), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n659), .B1(new_n797), .B2(KEYINPUT116), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n798), .A2(KEYINPUT117), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT117), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n794), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n706), .A2(new_n643), .A3(new_n657), .A4(new_n735), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n761), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n809), .A2(new_n634), .A3(new_n710), .ZN(new_n810));
  INV_X1    g624(.A(new_n234), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n675), .A2(new_n676), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n587), .A4(new_n612), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT51), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT51), .B1(new_n815), .B2(KEYINPUT118), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(KEYINPUT118), .B2(new_n815), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n806), .A3(new_n796), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n813), .A3(new_n613), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n745), .A2(new_n809), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT48), .Z(new_n823));
  INV_X1    g637(.A(G952), .ZN(new_n824));
  INV_X1    g638(.A(new_n716), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n824), .B(G953), .C1(new_n794), .C2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n821), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n817), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n657), .A2(new_n444), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n645), .A2(new_n590), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n667), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n734), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n675), .B2(new_n676), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n719), .B1(new_n641), .B2(new_n648), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n691), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n829), .B(KEYINPUT52), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n719), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n649), .A2(new_n691), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n734), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n357), .A2(new_n674), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT96), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n357), .A2(new_n670), .A3(new_n674), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n837), .B1(new_n840), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n836), .B2(new_n829), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n838), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n633), .A2(new_n537), .A3(new_n645), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n625), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n437), .A2(new_n754), .A3(new_n853), .A4(new_n590), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n851), .B1(new_n783), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n754), .A2(new_n853), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n641), .A2(KEYINPUT111), .A3(new_n595), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n718), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n737), .B2(new_n738), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n752), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n641), .B(new_n811), .C1(new_n696), .C2(new_n591), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n613), .B(KEYINPUT109), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n536), .A2(new_n587), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n493), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n599), .A3(new_n590), .A4(new_n437), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n713), .A2(new_n868), .A3(new_n636), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n862), .A2(new_n869), .A3(new_n701), .A4(new_n704), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n749), .A2(new_n861), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT52), .B1(new_n840), .B2(new_n845), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n834), .A2(new_n835), .A3(new_n848), .A4(new_n691), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n744), .B(new_n717), .C1(new_n738), .C2(new_n737), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n641), .A2(new_n811), .ZN(new_n877));
  INV_X1    g691(.A(new_n738), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n734), .A2(KEYINPUT102), .A3(new_n736), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI22_X1  g694(.A1(KEYINPUT42), .A2(new_n876), .B1(new_n880), .B2(new_n747), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n701), .A2(new_n862), .A3(new_n869), .A4(new_n704), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n752), .A2(new_n858), .A3(new_n860), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n885));
  AOI22_X1  g699(.A1(new_n850), .A2(new_n872), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n884), .A2(new_n885), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n749), .A2(new_n870), .A3(new_n861), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT112), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n883), .A3(new_n882), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n850), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n895), .B2(new_n871), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n888), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n792), .B1(new_n828), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n760), .A2(new_n234), .A3(new_n735), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT108), .Z(new_n900));
  AOI211_X1 g714(.A(new_n659), .B(new_n900), .C1(KEYINPUT49), .C2(new_n706), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n901), .B(new_n813), .C1(KEYINPUT49), .C2(new_n706), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n218), .A2(G952), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT120), .Z(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n886), .A2(new_n188), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n457), .A2(new_n473), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n471), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT55), .Z(new_n911));
  OR2_X1    g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n911), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(G51));
  NOR3_X1   g728(.A1(new_n886), .A2(new_n188), .A3(new_n774), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT121), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n847), .A2(new_n849), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n846), .A2(KEYINPUT113), .A3(new_n848), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n873), .A2(new_n874), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n885), .B1(new_n892), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n888), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n360), .B(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n435), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n904), .B1(new_n916), .B2(new_n927), .ZN(G54));
  NAND3_X1  g742(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n568), .A3(new_n580), .ZN(new_n930));
  INV_X1    g744(.A(new_n904), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n907), .A2(KEYINPUT58), .A3(G475), .A4(new_n581), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(G60));
  AND2_X1   g747(.A1(new_n608), .A2(new_n610), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n602), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n897), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n924), .A2(new_n935), .A3(new_n937), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n938), .A2(new_n939), .A3(new_n906), .ZN(G63));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n187), .A2(new_n188), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n922), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n944), .ZN(new_n946));
  AOI211_X1 g760(.A(KEYINPUT124), .B(new_n946), .C1(new_n919), .C2(new_n921), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n631), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT124), .B1(new_n886), .B2(new_n946), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n922), .A2(new_n941), .A3(new_n944), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n231), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n951), .A3(new_n905), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n948), .A2(new_n951), .A3(KEYINPUT61), .A4(new_n905), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  OAI21_X1  g770(.A(G953), .B1(new_n441), .B2(new_n466), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n882), .B2(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n909), .B1(G898), .B2(new_n218), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G69));
  NAND2_X1  g774(.A1(new_n328), .A2(new_n330), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n574), .A2(new_n575), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n840), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n679), .B2(new_n680), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n863), .A2(new_n866), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n877), .A2(new_n652), .A3(new_n755), .A4(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n789), .A2(new_n781), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n972), .B2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n881), .A2(new_n752), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n744), .A2(new_n715), .A3(new_n666), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n965), .B1(new_n780), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n789), .A2(new_n781), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n975), .A2(new_n218), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n218), .B1(G227), .B2(G900), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G72));
  NAND3_X1  g798(.A1(new_n975), .A2(new_n978), .A3(new_n882), .ZN(new_n985));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT126), .Z(new_n988));
  NAND2_X1  g802(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n326), .A3(new_n301), .A4(new_n331), .ZN(new_n990));
  INV_X1    g804(.A(new_n343), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n313), .B1(new_n331), .B2(new_n301), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n990), .B(new_n931), .C1(new_n896), .C2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n968), .A2(new_n971), .A3(new_n882), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n988), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n995), .B2(new_n988), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n997), .A2(new_n998), .A3(new_n671), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n994), .A2(new_n999), .ZN(G57));
endmodule


