

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  AND2_X1 U324 ( .A1(G229GAT), .A2(G233GAT), .ZN(n292) );
  NOR2_X1 U325 ( .A1(n543), .A2(n528), .ZN(n293) );
  XNOR2_X1 U326 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U327 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U328 ( .A(G113GAT), .B(G1GAT), .Z(n351) );
  XNOR2_X1 U329 ( .A(n422), .B(KEYINPUT54), .ZN(n423) );
  XNOR2_X1 U330 ( .A(n356), .B(n292), .ZN(n357) );
  XNOR2_X1 U331 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n403) );
  XNOR2_X1 U332 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U333 ( .A(n358), .B(n357), .ZN(n362) );
  XNOR2_X1 U334 ( .A(n404), .B(n403), .ZN(n535) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n463) );
  XNOR2_X1 U336 ( .A(n463), .B(KEYINPUT58), .ZN(n464) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT55), .B(KEYINPUT123), .Z(n444) );
  XOR2_X1 U339 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U340 ( .A(KEYINPUT95), .B(KEYINPUT1), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U342 ( .A(G85GAT), .B(G155GAT), .Z(n297) );
  XNOR2_X1 U343 ( .A(G29GAT), .B(G162GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U345 ( .A(G57GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n303) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U352 ( .A(KEYINPUT4), .B(n304), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n308) );
  XNOR2_X1 U355 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n431) );
  XOR2_X1 U357 ( .A(n309), .B(n431), .Z(n311) );
  XOR2_X1 U358 ( .A(G134GAT), .B(KEYINPUT0), .Z(n447) );
  XNOR2_X1 U359 ( .A(n351), .B(n447), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n550) );
  XOR2_X1 U362 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n315) );
  XNOR2_X1 U363 ( .A(KEYINPUT11), .B(KEYINPUT65), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U365 ( .A(n316), .B(KEYINPUT66), .Z(n318) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XNOR2_X1 U367 ( .A(G134GAT), .B(n438), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n324) );
  XOR2_X1 U369 ( .A(G92GAT), .B(G218GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(G190GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n408) );
  XOR2_X1 U372 ( .A(KEYINPUT9), .B(n408), .Z(n322) );
  NAND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(n324), .B(n323), .Z(n332) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n326) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(G29GAT), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U379 ( .A(KEYINPUT8), .B(n327), .Z(n366) );
  XOR2_X1 U380 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n329) );
  XNOR2_X1 U381 ( .A(G106GAT), .B(G85GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U383 ( .A(G99GAT), .B(n330), .Z(n373) );
  XNOR2_X1 U384 ( .A(n366), .B(n373), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n563) );
  XOR2_X1 U386 ( .A(KEYINPUT15), .B(G64GAT), .Z(n334) );
  XNOR2_X1 U387 ( .A(G211GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT13), .Z(n378) );
  XOR2_X1 U390 ( .A(n335), .B(n378), .Z(n337) );
  XNOR2_X1 U391 ( .A(G1GAT), .B(G71GAT), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n338), .B(KEYINPUT82), .ZN(n412) );
  XOR2_X1 U395 ( .A(n339), .B(n412), .Z(n341) );
  XOR2_X1 U396 ( .A(G15GAT), .B(G127GAT), .Z(n451) );
  XOR2_X1 U397 ( .A(G22GAT), .B(G155GAT), .Z(n437) );
  XNOR2_X1 U398 ( .A(n451), .B(n437), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U400 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n343) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U403 ( .A(n345), .B(n344), .Z(n350) );
  XOR2_X1 U404 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n347) );
  XNOR2_X1 U405 ( .A(KEYINPUT83), .B(KEYINPUT86), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n348), .B(KEYINPUT87), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n585) );
  NAND2_X1 U409 ( .A1(n563), .A2(n585), .ZN(n393) );
  XOR2_X1 U410 ( .A(G36GAT), .B(G50GAT), .Z(n353) );
  XNOR2_X1 U411 ( .A(n351), .B(KEYINPUT67), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U413 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n355) );
  XNOR2_X1 U414 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G141GAT), .Z(n360) );
  XNOR2_X1 U417 ( .A(G197GAT), .B(G22GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U419 ( .A(n362), .B(n361), .Z(n368) );
  XOR2_X1 U420 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n364) );
  XNOR2_X1 U421 ( .A(G169GAT), .B(G8GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n577) );
  XOR2_X1 U425 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XNOR2_X1 U426 ( .A(G176GAT), .B(G204GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n369), .B(G64GAT), .ZN(n411) );
  XOR2_X1 U428 ( .A(n448), .B(n411), .Z(n371) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n387) );
  XOR2_X1 U432 ( .A(KEYINPUT33), .B(KEYINPUT79), .Z(n375) );
  XNOR2_X1 U433 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n377) );
  INV_X1 U435 ( .A(KEYINPUT73), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n378), .B(G92GAT), .ZN(n379) );
  XNOR2_X1 U438 ( .A(n380), .B(n379), .ZN(n382) );
  INV_X1 U439 ( .A(KEYINPUT74), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n385) );
  XNOR2_X1 U441 ( .A(G78GAT), .B(KEYINPUT76), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n383), .B(G148GAT), .ZN(n435) );
  XNOR2_X1 U443 ( .A(n435), .B(KEYINPUT32), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n399) );
  XNOR2_X1 U446 ( .A(n399), .B(KEYINPUT41), .ZN(n570) );
  NOR2_X1 U447 ( .A1(n577), .A2(n570), .ZN(n391) );
  XNOR2_X1 U448 ( .A(KEYINPUT46), .B(KEYINPUT117), .ZN(n389) );
  INV_X1 U449 ( .A(KEYINPUT116), .ZN(n388) );
  NOR2_X1 U450 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U451 ( .A(KEYINPUT47), .B(n394), .ZN(n396) );
  INV_X1 U452 ( .A(KEYINPUT118), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n396), .B(n395), .ZN(n402) );
  XOR2_X1 U454 ( .A(KEYINPUT81), .B(n563), .Z(n543) );
  XNOR2_X1 U455 ( .A(KEYINPUT36), .B(n543), .ZN(n590) );
  NOR2_X1 U456 ( .A1(n585), .A2(n590), .ZN(n397) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(n397), .ZN(n398) );
  NAND2_X1 U458 ( .A1(n398), .A2(n577), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n400), .A2(n399), .ZN(n401) );
  NOR2_X1 U460 ( .A1(n402), .A2(n401), .ZN(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n406) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n420) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n418) );
  XOR2_X1 U468 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n414) );
  XNOR2_X1 U469 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n455) );
  XOR2_X1 U471 ( .A(G211GAT), .B(KEYINPUT21), .Z(n416) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(KEYINPUT91), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n432) );
  XNOR2_X1 U474 ( .A(n455), .B(n432), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n498) );
  XNOR2_X1 U477 ( .A(n498), .B(KEYINPUT121), .ZN(n421) );
  NOR2_X1 U478 ( .A1(n535), .A2(n421), .ZN(n424) );
  INV_X1 U479 ( .A(KEYINPUT122), .ZN(n422) );
  NOR2_X1 U480 ( .A1(n550), .A2(n425), .ZN(n576) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n427) );
  XNOR2_X1 U482 ( .A(G218GAT), .B(G106GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n442) );
  XOR2_X1 U484 ( .A(G204GAT), .B(KEYINPUT93), .Z(n429) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U487 ( .A(n430), .B(KEYINPUT24), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U490 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n470) );
  NAND2_X1 U494 ( .A1(n576), .A2(n470), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n566) );
  XOR2_X1 U496 ( .A(KEYINPUT90), .B(G190GAT), .Z(n446) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G99GAT), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n462) );
  XOR2_X1 U499 ( .A(n448), .B(n447), .Z(n450) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U502 ( .A(n452), .B(n451), .Z(n460) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G183GAT), .Z(n454) );
  XNOR2_X1 U504 ( .A(G113GAT), .B(KEYINPUT89), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT88), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n456), .B(KEYINPUT20), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U509 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U510 ( .A(n462), .B(n461), .ZN(n565) );
  INV_X1 U511 ( .A(n565), .ZN(n528) );
  AND2_X1 U512 ( .A1(n566), .A2(n293), .ZN(n465) );
  INV_X1 U513 ( .A(n550), .ZN(n521) );
  NOR2_X1 U514 ( .A1(n577), .A2(n399), .ZN(n493) );
  XOR2_X1 U515 ( .A(n498), .B(KEYINPUT27), .Z(n469) );
  XNOR2_X1 U516 ( .A(n470), .B(KEYINPUT28), .ZN(n532) );
  NAND2_X1 U517 ( .A1(n550), .A2(n532), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n469), .A2(n466), .ZN(n536) );
  NAND2_X1 U519 ( .A1(n528), .A2(n536), .ZN(n476) );
  NAND2_X1 U520 ( .A1(n498), .A2(n565), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n470), .A2(n467), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n468), .Z(n473) );
  INV_X1 U523 ( .A(n469), .ZN(n472) );
  NOR2_X1 U524 ( .A1(n565), .A2(n470), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT26), .ZN(n575) );
  NAND2_X1 U526 ( .A1(n472), .A2(n575), .ZN(n548) );
  NAND2_X1 U527 ( .A1(n473), .A2(n548), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n521), .A2(n474), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n476), .A2(n475), .ZN(n489) );
  INV_X1 U530 ( .A(n585), .ZN(n559) );
  NAND2_X1 U531 ( .A1(n543), .A2(n559), .ZN(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U533 ( .A1(n489), .A2(n478), .ZN(n507) );
  NAND2_X1 U534 ( .A1(n493), .A2(n507), .ZN(n486) );
  NOR2_X1 U535 ( .A1(n521), .A2(n486), .ZN(n480) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  INV_X1 U539 ( .A(n498), .ZN(n525) );
  NOR2_X1 U540 ( .A1(n525), .A2(n486), .ZN(n482) );
  XOR2_X1 U541 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U542 ( .A1(n528), .A2(n486), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n532), .A2(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n496) );
  NAND2_X1 U550 ( .A1(n585), .A2(n489), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(n490), .ZN(n491) );
  NOR2_X1 U552 ( .A1(n590), .A2(n491), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n492), .Z(n520) );
  NAND2_X1 U554 ( .A1(n520), .A2(n493), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(n494), .Z(n502) );
  NAND2_X1 U556 ( .A1(n502), .A2(n550), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U558 ( .A(G29GAT), .B(n497), .Z(G1328GAT) );
  NAND2_X1 U559 ( .A1(n502), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n502), .A2(n565), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT40), .ZN(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n505) );
  INV_X1 U565 ( .A(n532), .ZN(n503) );
  NAND2_X1 U566 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  INV_X1 U569 ( .A(n577), .ZN(n552) );
  NOR2_X1 U570 ( .A1(n552), .A2(n570), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n519), .A2(n507), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n521), .A2(n514), .ZN(n509) );
  XNOR2_X1 U573 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n510), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n525), .A2(n514), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n528), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n532), .ZN(n518) );
  XOR2_X1 U582 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n516) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT111), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NAND2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n531) );
  NOR2_X1 U587 ( .A1(n521), .A2(n531), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n531), .ZN(n526) );
  XOR2_X1 U592 ( .A(KEYINPUT114), .B(n526), .Z(n527) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n531), .ZN(n530) );
  XNOR2_X1 U595 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n536), .A2(n565), .ZN(n537) );
  NOR2_X1 U601 ( .A1(n535), .A2(n537), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n552), .A2(n545), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  INV_X1 U605 ( .A(n570), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n545), .A2(n555), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n559), .A2(n545), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  INV_X1 U612 ( .A(n543), .ZN(n544) );
  NAND2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n535), .A2(n548), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT119), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n552), .A2(n561), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U627 ( .A(n561), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n573) );
  NOR2_X1 U631 ( .A1(n577), .A2(n573), .ZN(n567) );
  XOR2_X1 U632 ( .A(G169GAT), .B(n567), .Z(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n572) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1349GAT) );
  NOR2_X1 U638 ( .A1(n585), .A2(n573), .ZN(n574) );
  XOR2_X1 U639 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n589) );
  NOR2_X1 U641 ( .A1(n589), .A2(n577), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n589), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n582), .A2(n399), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n589), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

