//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  XNOR2_X1  g000(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(G143), .A4(G214), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT18), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(G131), .ZN(new_n204));
  OAI221_X1 g018(.A(new_n193), .B1(new_n200), .B2(new_n203), .C1(new_n204), .C2(new_n201), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT16), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT71), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT71), .A4(KEYINPUT16), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(G146), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT72), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n213), .A2(new_n214), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G146), .A4(new_n212), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n214), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT71), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n192), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n200), .A2(KEYINPUT17), .A3(G131), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n216), .A2(new_n219), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT86), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n200), .B2(G131), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n198), .A2(KEYINPUT86), .A3(new_n202), .A4(new_n199), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n204), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n224), .B2(new_n225), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n190), .B(new_n205), .C1(new_n226), .C2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n191), .B(KEYINPUT19), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n192), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(new_n204), .A3(new_n230), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n215), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n205), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n190), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(G475), .A2(G902), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n187), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  AOI211_X1 g060(.A(KEYINPUT20), .B(new_n246), .C1(new_n233), .C2(new_n242), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n205), .B1(new_n226), .B2(new_n232), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n241), .ZN(new_n249));
  AOI21_X1  g063(.A(G902), .B1(new_n249), .B2(new_n233), .ZN(new_n250));
  INV_X1    g064(.A(G475), .ZN(new_n251));
  OAI22_X1  g065(.A1(new_n245), .A2(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT89), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n254));
  OAI221_X1 g068(.A(new_n254), .B1(new_n250), .B2(new_n251), .C1(new_n245), .C2(new_n247), .ZN(new_n255));
  INV_X1    g069(.A(G902), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  INV_X1    g071(.A(G122), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G116), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n259), .B2(KEYINPUT14), .ZN(new_n260));
  INV_X1    g074(.A(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G122), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n260), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT66), .B(G128), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n197), .A2(G128), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n268), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G134), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n264), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT13), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n265), .A2(G143), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT90), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n197), .A2(KEYINPUT13), .A3(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n274), .A2(KEYINPUT90), .ZN(new_n278));
  OAI21_X1  g092(.A(G134), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n263), .A2(new_n257), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n259), .A2(new_n262), .A3(G107), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n272), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT9), .B(G234), .ZN(new_n285));
  INV_X1    g099(.A(G217), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n285), .A2(new_n286), .A3(G953), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n274), .A2(KEYINPUT90), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n275), .A3(new_n276), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n282), .B1(new_n290), .B2(G134), .ZN(new_n291));
  INV_X1    g105(.A(new_n287), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n272), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n256), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G478), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(KEYINPUT15), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n292), .B1(new_n291), .B2(new_n272), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n284), .A2(new_n287), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n296), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n256), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(KEYINPUT91), .A2(G952), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT91), .A2(G952), .ZN(new_n306));
  AOI21_X1  g120(.A(G953), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G234), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(new_n194), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n256), .B(new_n195), .C1(G234), .C2(G237), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT21), .B(G898), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n303), .A2(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n253), .A2(new_n255), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n316), .B(KEYINPUT79), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G210), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n320));
  INV_X1    g134(.A(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G116), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n261), .A2(G119), .ZN(new_n323));
  INV_X1    g137(.A(G113), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n322), .B(new_n323), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(new_n323), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n257), .A3(G104), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n189), .A2(G107), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G101), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n336), .A2(G101), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n332), .A2(new_n334), .A3(new_n340), .A4(new_n335), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n331), .B(new_n338), .C1(new_n339), .C2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT5), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(G113), .C1(KEYINPUT5), .C2(new_n322), .ZN(new_n345));
  INV_X1    g159(.A(new_n335), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n189), .A2(G107), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n327), .A3(new_n348), .A4(new_n341), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G122), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(KEYINPUT80), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n353), .B1(new_n343), .B2(new_n349), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT82), .A3(new_n351), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n343), .A2(new_n349), .A3(new_n352), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n361));
  OAI211_X1 g175(.A(KEYINPUT6), .B(new_n360), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(KEYINPUT81), .B(new_n353), .C1(new_n343), .C2(new_n349), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n357), .B(new_n359), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n192), .A2(G143), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n197), .A2(G146), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(KEYINPUT0), .A2(G128), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT0), .ZN(new_n369));
  INV_X1    g183(.A(G128), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G143), .B(G146), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n369), .B2(new_n370), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G125), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(G143), .B2(new_n192), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n367), .B1(new_n265), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n370), .A2(KEYINPUT1), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n365), .A3(new_n366), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n376), .B1(new_n383), .B2(G125), .ZN(new_n384));
  INV_X1    g198(.A(G224), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n384), .B(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n320), .B1(new_n364), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n359), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT82), .B1(new_n358), .B2(new_n351), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n350), .A2(new_n354), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n358), .A2(new_n361), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n394), .A4(new_n360), .ZN(new_n395));
  INV_X1    g209(.A(new_n387), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT83), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n386), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n384), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n399), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n345), .A2(new_n327), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n348), .A2(new_n341), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n349), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n352), .B(KEYINPUT8), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n401), .A2(new_n360), .A3(new_n402), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n256), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n319), .B1(new_n398), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n319), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n413), .B(new_n410), .C1(new_n388), .C2(new_n397), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n318), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G221), .B1(new_n285), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT76), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n381), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n380), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G128), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n423), .B1(new_n367), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT77), .B1(new_n426), .B2(new_n404), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n367), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT76), .B1(new_n373), .B2(new_n380), .ZN(new_n429));
  AND4_X1   g243(.A1(KEYINPUT76), .A2(new_n380), .A3(new_n365), .A4(new_n366), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n404), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT10), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G137), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT64), .B1(new_n436), .B2(G134), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n267), .B2(G137), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n267), .A3(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(KEYINPUT11), .A3(G134), .ZN(new_n442));
  AND4_X1   g256(.A1(new_n437), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n202), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n437), .A2(new_n439), .A3(new_n441), .A4(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G131), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT10), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n379), .B2(new_n381), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n432), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n339), .A2(new_n342), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n375), .A2(new_n338), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n435), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n426), .A2(KEYINPUT77), .A3(new_n404), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n456));
  OAI22_X1  g270(.A1(new_n455), .A2(new_n456), .B1(new_n382), .B2(new_n432), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT12), .A3(new_n447), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n427), .A2(new_n434), .B1(new_n383), .B2(new_n404), .ZN(new_n460));
  INV_X1    g274(.A(new_n447), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n454), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT75), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n195), .A2(G227), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n468));
  INV_X1    g282(.A(new_n453), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT78), .B1(new_n435), .B2(new_n453), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n469), .A3(new_n461), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n463), .A2(new_n467), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n420), .B1(new_n476), .B2(new_n256), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n467), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n473), .B2(new_n454), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n458), .A2(new_n462), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n474), .A3(new_n467), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n420), .A3(new_n256), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n419), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT84), .B(new_n318), .C1(new_n412), .C2(new_n414), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n315), .A2(new_n417), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n194), .A2(new_n195), .A3(G210), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT27), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT26), .B(G101), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n444), .A2(new_n446), .B1(new_n372), .B2(new_n374), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n267), .A2(KEYINPUT65), .A3(G137), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT65), .B1(new_n267), .B2(G137), .ZN(new_n494));
  OAI22_X1  g308(.A1(new_n493), .A2(new_n494), .B1(new_n267), .B2(G137), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G131), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n202), .A2(new_n443), .B1(new_n379), .B2(new_n381), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n492), .A2(KEYINPUT67), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n331), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n445), .A2(G131), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n445), .A2(G131), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n375), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n444), .A2(new_n382), .A3(new_n496), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n502), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n447), .A2(KEYINPUT67), .A3(new_n375), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n509), .A3(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n508), .B1(new_n510), .B2(KEYINPUT30), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n491), .B(new_n505), .C1(new_n511), .C2(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n506), .B1(new_n498), .B2(new_n504), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n331), .B1(new_n514), .B2(new_n508), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n491), .A4(new_n505), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(KEYINPUT31), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n502), .A2(new_n507), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n505), .B1(new_n499), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n499), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n491), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n512), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G472), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n256), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT32), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n530), .A2(new_n534), .A3(new_n531), .A4(new_n256), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n515), .A2(new_n505), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n526), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n537), .B(new_n538), .C1(new_n526), .C2(new_n525), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n510), .A2(new_n331), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n505), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n541), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(KEYINPUT28), .B1(KEYINPUT70), .B2(new_n524), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n491), .A2(KEYINPUT29), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n539), .B(new_n256), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n533), .A2(new_n535), .B1(G472), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n191), .A2(new_n192), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n370), .A2(G119), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n265), .B2(G119), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT24), .B(G110), .Z(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n265), .A2(KEYINPUT23), .A3(G119), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT23), .B1(new_n370), .B2(G119), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n321), .B2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n552), .A2(KEYINPUT73), .B1(new_n556), .B2(G110), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n215), .B(new_n548), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n216), .A2(new_n219), .A3(new_n222), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n556), .A2(G110), .B1(new_n550), .B2(new_n551), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT74), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n567), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n286), .B1(G234), .B2(new_n256), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n568), .A2(new_n576), .A3(new_n256), .A4(new_n570), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT25), .B1(new_n571), .B2(G902), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OR3_X1    g395(.A1(new_n487), .A2(new_n547), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  NAND2_X1  g397(.A1(new_n530), .A2(new_n256), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G472), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n532), .A3(new_n485), .A4(new_n580), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT92), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n253), .A2(new_n255), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n300), .A2(new_n295), .A3(new_n256), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n298), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n592), .A2(new_n300), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n300), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n589), .B1(new_n595), .B2(new_n295), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n313), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n599), .B(new_n318), .C1(new_n412), .C2(new_n414), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n587), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT94), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NAND2_X1  g419(.A1(new_n398), .A2(new_n411), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n413), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n398), .A2(new_n319), .A3(new_n411), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n317), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n246), .B1(new_n233), .B2(new_n242), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n187), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT95), .B1(new_n610), .B2(new_n187), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n303), .B1(new_n250), .B2(new_n251), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n610), .A2(new_n616), .A3(new_n187), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n609), .A2(new_n618), .A3(new_n619), .A4(new_n599), .ZN(new_n620));
  INV_X1    g434(.A(new_n615), .ZN(new_n621));
  INV_X1    g435(.A(new_n617), .ZN(new_n622));
  INV_X1    g436(.A(new_n245), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(KEYINPUT95), .A3(new_n611), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT96), .B1(new_n600), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n587), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NAND2_X1  g444(.A1(new_n578), .A2(new_n579), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n563), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n573), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n585), .A2(new_n532), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n487), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT37), .B(G110), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n609), .A2(new_n635), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n533), .A2(new_n535), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n546), .A2(G472), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n310), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n309), .B1(G900), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT97), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n643), .A2(new_n485), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n513), .A2(new_n517), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n526), .B2(new_n541), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n651), .B2(G902), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n646), .B(KEYINPUT39), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n485), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT40), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n412), .A2(new_n414), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n635), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n318), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n588), .A2(new_n303), .ZN(new_n663));
  OR4_X1    g477(.A1(new_n654), .A2(new_n657), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(new_n646), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n588), .A2(new_n597), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n596), .B1(new_n253), .B2(new_n255), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(KEYINPUT99), .A3(new_n666), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n643), .A2(new_n485), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NAND2_X1  g487(.A1(new_n641), .A2(new_n642), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n470), .B1(new_n468), .B2(new_n469), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n453), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n447), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n467), .B1(new_n677), .B2(new_n474), .ZN(new_n678));
  INV_X1    g492(.A(new_n482), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n256), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n420), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n483), .B(new_n256), .C1(new_n681), .C2(new_n420), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n683), .A2(new_n684), .A3(new_n418), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n601), .A3(new_n580), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND4_X1  g502(.A1(new_n627), .A2(new_n674), .A3(new_n580), .A4(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NAND3_X1  g504(.A1(new_n685), .A2(KEYINPUT101), .A3(new_n609), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n683), .A2(new_n684), .A3(new_n418), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n692), .B1(new_n693), .B2(new_n415), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n661), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n253), .A2(new_n255), .A3(new_n314), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n641), .B2(new_n642), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT103), .B(G119), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G21));
  NOR2_X1   g518(.A1(new_n663), .A2(new_n415), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n526), .B1(new_n542), .B2(new_n543), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n518), .A2(new_n706), .A3(new_n529), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n707), .A2(new_n531), .A3(new_n256), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n531), .B1(new_n530), .B2(new_n256), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n581), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n705), .A2(new_n599), .A3(new_n685), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n695), .A2(new_n669), .A3(new_n671), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n485), .A2(new_n318), .A3(new_n658), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n674), .A2(new_n718), .A3(new_n580), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n669), .A2(new_n671), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n547), .A2(new_n581), .A3(new_n717), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n667), .A2(new_n668), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT99), .B1(new_n670), .B2(new_n666), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n725), .A3(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  XNOR2_X1  g542(.A(new_n647), .B(KEYINPUT104), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT105), .B(G134), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G36));
  NAND2_X1  g546(.A1(new_n658), .A2(new_n318), .ZN(new_n733));
  INV_X1    g547(.A(new_n588), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n597), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n661), .B1(new_n585), .B2(new_n532), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n733), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n739), .A2(KEYINPUT44), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n744), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n476), .B(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(G469), .ZN(new_n750));
  NAND2_X1  g564(.A1(G469), .A2(G902), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n749), .C2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n484), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(new_n418), .A3(new_n655), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n747), .A2(new_n748), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT107), .B(G137), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G39));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n418), .ZN(new_n760));
  XOR2_X1   g574(.A(new_n760), .B(KEYINPUT47), .Z(new_n761));
  NOR3_X1   g575(.A1(new_n674), .A2(new_n580), .A3(new_n733), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n725), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  NOR4_X1   g578(.A1(new_n660), .A2(new_n581), .A3(new_n419), .A4(new_n317), .ZN(new_n765));
  INV_X1    g579(.A(new_n735), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n683), .A2(new_n684), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT49), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n654), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n738), .A2(new_n309), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n710), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n691), .A2(new_n694), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n733), .A2(new_n693), .A3(new_n581), .A4(new_n309), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n654), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT114), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n773), .B(new_n307), .C1(new_n598), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n547), .A2(new_n581), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n733), .A2(new_n693), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n770), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT48), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(KEYINPUT48), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT117), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n777), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n733), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n767), .A2(new_n419), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n771), .B(new_n787), .C1(new_n761), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(KEYINPUT51), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n660), .A2(new_n318), .A3(new_n693), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n770), .A2(new_n710), .A3(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT113), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n771), .A2(KEYINPUT50), .A3(new_n791), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n708), .A2(new_n709), .A3(new_n661), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n770), .A2(new_n800), .A3(new_n779), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n734), .A2(new_n596), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n776), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n790), .A2(new_n799), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n799), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n789), .B(new_n801), .C1(new_n776), .C2(new_n802), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n786), .B(new_n806), .C1(new_n809), .C2(KEYINPUT51), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n695), .A2(new_n697), .A3(new_n700), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n700), .B1(new_n695), .B2(new_n697), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n689), .A2(new_n686), .A3(new_n711), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT108), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n417), .A2(new_n599), .A3(new_n486), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n253), .A2(new_n255), .A3(new_n303), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n817), .A2(new_n586), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT110), .B1(new_n819), .B2(new_n637), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n417), .A2(new_n486), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n599), .A4(new_n670), .ZN(new_n823));
  INV_X1    g637(.A(new_n532), .ZN(new_n824));
  AOI211_X1 g638(.A(G469), .B(G902), .C1(new_n480), .C2(new_n482), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n580), .B(new_n418), .C1(new_n825), .C2(new_n477), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n824), .A2(new_n826), .A3(new_n709), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT109), .B1(new_n817), .B2(new_n598), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n636), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n821), .A2(new_n830), .A3(new_n315), .A4(new_n485), .ZN(new_n831));
  INV_X1    g645(.A(new_n818), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n821), .A2(new_n599), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n582), .A2(new_n820), .A3(new_n829), .A4(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n689), .A2(new_n686), .A3(new_n711), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT108), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n702), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n816), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n303), .A2(new_n646), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n251), .B2(new_n250), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n842), .A2(new_n661), .A3(new_n617), .A4(new_n614), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n674), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n800), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n844), .B1(new_n720), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n846), .A2(new_n718), .B1(new_n722), .B2(new_n729), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n727), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n631), .A2(new_n634), .A3(new_n666), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT111), .Z(new_n850));
  NAND4_X1  g664(.A1(new_n653), .A2(new_n705), .A3(new_n485), .A4(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n714), .A2(new_n672), .A3(new_n648), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n485), .B(new_n643), .C1(new_n725), .C2(new_n647), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n714), .A4(new_n851), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n848), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n856), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n847), .A2(new_n727), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n816), .A2(new_n836), .A3(new_n839), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n811), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n727), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n820), .A2(new_n835), .A3(new_n829), .A4(new_n582), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n866), .A2(new_n867), .A3(new_n859), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n847), .A2(new_n702), .A3(new_n837), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n860), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n864), .A2(new_n811), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n810), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT118), .Z(new_n874));
  OAI21_X1  g688(.A(new_n769), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT119), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n877), .B(new_n769), .C1(new_n872), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(G75));
  NAND2_X1  g693(.A1(new_n864), .A2(new_n870), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(G210), .A3(G902), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n387), .B(KEYINPUT55), .Z(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n364), .B(KEYINPUT120), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT121), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n886), .B2(new_n887), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n195), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  XOR2_X1   g707(.A(new_n751), .B(KEYINPUT57), .Z(new_n894));
  AOI21_X1  g708(.A(new_n811), .B1(new_n864), .B2(new_n870), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n871), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n483), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n880), .A2(G902), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n898), .A2(new_n750), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n892), .B1(new_n897), .B2(new_n899), .ZN(G54));
  INV_X1    g714(.A(new_n892), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n898), .A2(new_n902), .A3(new_n251), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n903), .B2(new_n243), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n243), .B2(new_n903), .ZN(G60));
  NAND2_X1  g719(.A1(new_n593), .A2(new_n594), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n871), .A2(new_n865), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n840), .B2(new_n857), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n868), .A2(new_n860), .A3(new_n869), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n864), .A2(new_n811), .A3(new_n870), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n892), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n912), .B1(new_n871), .B2(new_n895), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n901), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT123), .B(new_n911), .C1(new_n919), .C2(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G63));
  INV_X1    g741(.A(new_n880), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n633), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n571), .B1(new_n928), .B2(new_n930), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n901), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g749(.A(G953), .B1(new_n311), .B2(new_n385), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n840), .B2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n888), .B1(G898), .B2(new_n195), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  AND2_X1   g754(.A1(new_n855), .A2(new_n714), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n756), .A2(new_n778), .A3(new_n705), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n763), .A2(new_n730), .A3(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(new_n727), .A2(new_n757), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n195), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n234), .B(KEYINPUT125), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n511), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(G900), .A2(G953), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n941), .A2(new_n664), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  INV_X1    g765(.A(new_n763), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n733), .B(new_n656), .C1(new_n598), .C2(new_n818), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n778), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n757), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n951), .A2(new_n757), .A3(KEYINPUT126), .A4(new_n954), .ZN(new_n958));
  AOI21_X1  g772(.A(G953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n949), .B1(new_n959), .B2(new_n947), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n949), .B(new_n963), .C1(new_n959), .C2(new_n947), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G72));
  INV_X1    g779(.A(new_n536), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n957), .A2(new_n840), .A3(new_n958), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT127), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n526), .B(new_n966), .C1(new_n967), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n537), .A2(new_n513), .A3(new_n517), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n969), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n858), .B2(new_n864), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n944), .B2(new_n840), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n966), .A2(new_n526), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n901), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n972), .A2(new_n975), .A3(new_n978), .ZN(G57));
endmodule


