//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n214));
  XOR2_X1   g0014(.A(new_n213), .B(new_n214), .Z(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  AND2_X1   g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n215), .A2(new_n228), .A3(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT8), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT66), .ZN(new_n257));
  OR3_X1    g0057(.A1(new_n222), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n209), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n253), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n251), .A2(new_n252), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n208), .B2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n269), .B2(G50), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT67), .ZN(new_n272));
  INV_X1    g0072(.A(new_n267), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n253), .B1(G1), .B2(new_n209), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n202), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n272), .B1(new_n264), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(new_n276), .A3(KEYINPUT9), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(new_n276), .A3(KEYINPUT68), .A4(KEYINPUT9), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G77), .ZN(new_n288));
  OAI211_X1 g0088(.A(G223), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n284), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n252), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  INV_X1    g0093(.A(G45), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(G1), .A3(G13), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n297), .A3(G274), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n217), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n292), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(G200), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n290), .B2(new_n291), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT69), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(G190), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n271), .A2(new_n276), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(KEYINPUT9), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n281), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n304), .B1(new_n303), .B2(G200), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n306), .A2(KEYINPUT69), .A3(new_n307), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT9), .B1(new_n271), .B2(new_n276), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n279), .A2(new_n280), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n209), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n329), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n222), .A2(new_n325), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n262), .A2(G159), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n324), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n287), .B2(new_n209), .ZN(new_n340));
  INV_X1    g0140(.A(new_n333), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n338), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n268), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n257), .A2(new_n258), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n274), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n266), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(G226), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n351));
  OAI211_X1 g0151(.A(G223), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n352));
  AND3_X1   g0152(.A1(KEYINPUT70), .A2(G33), .A3(G87), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT70), .B1(G33), .B2(G87), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n291), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT71), .B1(new_n356), .B2(new_n291), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n298), .B(new_n359), .C1(new_n223), .C2(new_n300), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n356), .A2(new_n291), .ZN(new_n362));
  INV_X1    g0162(.A(new_n300), .ZN(new_n363));
  INV_X1    g0163(.A(G274), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n231), .B2(new_n296), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n363), .A2(G232), .B1(new_n295), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(G200), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n345), .B(new_n350), .C1(new_n361), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT17), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n350), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n332), .A2(new_n333), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n338), .B1(new_n372), .B2(G68), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n253), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n374), .B2(new_n339), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n291), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n366), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n362), .A2(new_n366), .ZN(new_n381));
  INV_X1    g0181(.A(G169), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT18), .B1(new_n375), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n345), .A2(new_n350), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n357), .A2(new_n358), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n366), .A2(new_n378), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n382), .B2(new_n381), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n381), .A2(new_n307), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n377), .A2(new_n379), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n360), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n370), .A2(new_n385), .A3(new_n391), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G244), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n298), .B1(new_n397), .B2(new_n300), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n400));
  INV_X1    g0200(.A(G107), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n399), .B(new_n400), .C1(new_n401), .C2(new_n282), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(new_n291), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n378), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n255), .A2(new_n256), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n260), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n253), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n266), .ZN(new_n411));
  INV_X1    g0211(.A(G77), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n274), .B2(new_n412), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n404), .B1(G169), .B2(new_n403), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n403), .A2(G190), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n410), .A2(new_n414), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n307), .C2(new_n403), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n303), .A2(new_n382), .B1(new_n265), .B2(new_n270), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n306), .A2(new_n378), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n415), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n262), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n423), .A2(new_n202), .B1(new_n209), .B2(G68), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n259), .A2(new_n412), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n268), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT11), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT12), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n411), .B2(new_n325), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n274), .A2(new_n325), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n427), .B2(new_n426), .ZN(new_n434));
  OAI211_X1 g0234(.A(G232), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n435));
  OAI211_X1 g0235(.A(G226), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n291), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n363), .A2(G238), .B1(new_n295), .B2(new_n365), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(G179), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n443), .B1(new_n439), .B2(new_n440), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n445), .B1(new_n448), .B2(KEYINPUT14), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT14), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(new_n444), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(G169), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n434), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n451), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n434), .B1(new_n454), .B2(G190), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(G200), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n422), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NOR3_X1   g0258(.A1(new_n323), .A2(new_n396), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n208), .A2(G45), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n365), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n294), .A2(G1), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n297), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n469), .B2(new_n219), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(G264), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n472));
  OAI211_X1 g0272(.A(G257), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n473));
  INV_X1    g0273(.A(G303), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n282), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n475), .A2(new_n476), .A3(new_n291), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n475), .B2(new_n291), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n411), .A2(new_n218), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n208), .A2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n266), .A2(new_n481), .A3(new_n252), .A4(new_n251), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n482), .B2(new_n218), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT20), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n209), .B1(new_n224), .B2(G33), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT74), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G33), .A3(G283), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT74), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n218), .A2(G20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n268), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n484), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n487), .ZN(new_n494));
  INV_X1    g0294(.A(new_n485), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n268), .A2(new_n491), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT20), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n483), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT80), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n501), .B(new_n483), .C1(new_n493), .C2(new_n498), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n479), .B(G169), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT21), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n499), .B(KEYINPUT80), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(KEYINPUT21), .A3(G169), .A4(new_n479), .ZN(new_n507));
  OAI211_X1 g0307(.A(G179), .B(new_n471), .C1(new_n477), .C2(new_n478), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n500), .A2(new_n502), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n479), .A2(G200), .ZN(new_n512));
  OAI211_X1 g0312(.A(G190), .B(new_n471), .C1(new_n477), .C2(new_n478), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n505), .A2(new_n507), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n411), .A2(new_n224), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n482), .B2(new_n224), .ZN(new_n517));
  OAI21_X1  g0317(.A(G107), .B1(new_n340), .B2(new_n341), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT73), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT72), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n423), .A2(new_n412), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n401), .A2(KEYINPUT6), .A3(G97), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n521), .B(new_n523), .C1(new_n528), .C2(new_n209), .ZN(new_n529));
  AND2_X1   g0329(.A1(G97), .A2(G107), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n530), .B2(new_n205), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n209), .B1(new_n531), .B2(new_n524), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT72), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n372), .A2(KEYINPUT73), .A3(G107), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n520), .A2(new_n529), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n517), .B1(new_n535), .B2(new_n268), .ZN(new_n536));
  OAI211_X1 g0336(.A(G244), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G250), .A2(G1698), .ZN(new_n540));
  NAND2_X1  g0340(.A1(KEYINPUT4), .A2(G244), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n282), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n494), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n291), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT75), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n461), .A2(new_n462), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n291), .B1(new_n465), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(G257), .B1(new_n365), .B2(new_n463), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n537), .A2(new_n538), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n282), .A2(new_n542), .B1(new_n487), .B2(new_n489), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n297), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n464), .B1(new_n469), .B2(new_n225), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT75), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n555), .A3(G190), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n536), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n535), .A2(new_n268), .ZN(new_n560));
  INV_X1    g0360(.A(new_n517), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT76), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n546), .B1(new_n545), .B2(new_n549), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT75), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n382), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n553), .A2(new_n554), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n378), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n536), .A2(KEYINPUT76), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n559), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n297), .A2(G274), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n572), .B1(new_n573), .B2(new_n460), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n465), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n397), .A2(G1698), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(G238), .B2(G1698), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n578), .A2(new_n287), .B1(new_n327), .B2(new_n218), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n291), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n297), .A2(G250), .A3(new_n460), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n576), .A2(new_n580), .A3(G190), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT78), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n327), .A2(new_n218), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G238), .A2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n397), .B2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n585), .B1(new_n587), .B2(new_n282), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n581), .B1(new_n588), .B2(new_n297), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT77), .B1(new_n365), .B2(new_n465), .ZN(new_n590));
  AND4_X1   g0390(.A1(KEYINPUT77), .A2(new_n297), .A3(G274), .A4(new_n465), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n209), .B1(new_n437), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G87), .B2(new_n206), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n209), .B(G68), .C1(new_n285), .C2(new_n286), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n594), .B1(new_n259), .B2(new_n224), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n268), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n407), .A2(new_n411), .ZN(new_n601));
  INV_X1    g0401(.A(G87), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n482), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n581), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n579), .B2(new_n291), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT78), .A3(new_n576), .A4(G190), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n584), .A2(new_n593), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n606), .A2(new_n576), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n382), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n600), .B(new_n601), .C1(new_n407), .C2(new_n482), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n606), .A2(new_n378), .A3(new_n576), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n616));
  OAI211_X1 g0416(.A(G250), .B(new_n283), .C1(new_n285), .C2(new_n286), .ZN(new_n617));
  INV_X1    g0417(.A(G294), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n617), .C1(new_n327), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n291), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n548), .A2(G264), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n464), .A3(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(new_n378), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n619), .A2(new_n291), .B1(new_n548), .B2(G264), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n382), .B1(new_n624), .B2(new_n464), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n615), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n209), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n627));
  AND2_X1   g0427(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n628));
  NOR2_X1   g0428(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n282), .A2(new_n209), .A3(G87), .A4(new_n628), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT23), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n209), .B2(G107), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n401), .A2(KEYINPUT23), .A3(G20), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n634), .A2(new_n635), .B1(new_n585), .B2(new_n209), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT24), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT24), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n631), .A2(new_n632), .A3(new_n636), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n253), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n411), .A2(KEYINPUT25), .A3(new_n401), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT25), .B1(new_n411), .B2(new_n401), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(new_n401), .B2(new_n482), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n622), .A2(G169), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n624), .A2(G179), .A3(new_n464), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(KEYINPUT82), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n626), .A2(new_n645), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n641), .A2(new_n644), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n622), .A2(new_n307), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n624), .A2(new_n359), .A3(new_n464), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n614), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n459), .A2(new_n515), .A3(new_n571), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT83), .ZN(G372));
  NAND2_X1  g0457(.A1(new_n385), .A2(new_n391), .ZN(new_n658));
  INV_X1    g0458(.A(new_n457), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n453), .B1(new_n659), .B2(new_n415), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n370), .A2(new_n395), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n421), .B1(new_n663), .B2(new_n323), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n646), .A2(new_n647), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n645), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n507), .A2(new_n505), .A3(new_n510), .A4(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT84), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n604), .A2(new_n669), .A3(new_n593), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n307), .B1(new_n606), .B2(new_n576), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT84), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n673), .A3(new_n582), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n674), .A2(new_n654), .A3(new_n613), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT76), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n401), .B1(new_n332), .B2(new_n333), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(new_n519), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n529), .A2(new_n533), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n253), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n680), .B2(new_n517), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n550), .A2(new_n555), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n682), .A2(new_n382), .B1(new_n378), .B2(new_n566), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n570), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n668), .A2(new_n675), .A3(new_n684), .A4(new_n558), .ZN(new_n685));
  INV_X1    g0485(.A(new_n614), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT26), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n674), .A2(new_n613), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n536), .B1(new_n568), .B2(KEYINPUT85), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT85), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n688), .A2(new_n689), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n685), .A2(new_n613), .A3(new_n687), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n459), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n665), .A2(new_n695), .ZN(G369));
  AND2_X1   g0496(.A1(new_n507), .A2(new_n510), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n505), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n511), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g0507(.A(new_n515), .B(new_n698), .S(new_n707), .Z(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n649), .B(new_n654), .C1(new_n650), .C2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT86), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n649), .A2(new_n706), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n705), .B1(new_n697), .B2(new_n505), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n645), .A2(new_n666), .A3(new_n706), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n714), .A2(new_n718), .ZN(G399));
  NAND2_X1  g0519(.A1(new_n212), .A2(new_n293), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n230), .B2(new_n720), .ZN(new_n723));
  XOR2_X1   g0523(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n724));
  XNOR2_X1  g0524(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n613), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n684), .A2(new_n675), .A3(new_n558), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n697), .A2(new_n505), .A3(new_n649), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n690), .B1(new_n684), .B2(new_n686), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT26), .A4(new_n692), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n705), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n694), .A2(new_n706), .ZN(new_n734));
  XOR2_X1   g0534(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n735));
  AOI22_X1  g0535(.A1(new_n733), .A2(KEYINPUT29), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n589), .A2(new_n592), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n550), .A2(new_n555), .A3(new_n738), .A4(new_n624), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n508), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n739), .A2(new_n508), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT30), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n475), .A2(new_n291), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT79), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n475), .A2(new_n476), .A3(new_n291), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n470), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n609), .A2(new_n378), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n479), .A2(KEYINPUT90), .A3(new_n378), .A4(new_n609), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n566), .B1(new_n464), .B2(new_n624), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(KEYINPUT92), .B(new_n737), .C1(new_n739), .C2(new_n508), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n742), .A2(new_n744), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n705), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n571), .A2(new_n515), .A3(new_n655), .A4(new_n706), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n744), .A2(new_n754), .A3(new_n740), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n761), .A2(KEYINPUT91), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n763), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT91), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n759), .A2(new_n760), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n736), .B1(G330), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n725), .B1(new_n769), .B2(G1), .ZN(G364));
  INV_X1    g0570(.A(new_n720), .ZN(new_n771));
  INV_X1    g0571(.A(G13), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n208), .B1(new_n773), .B2(G45), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n708), .B2(G330), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G330), .B2(new_n708), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n212), .A2(new_n282), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(G116), .B2(new_n212), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n246), .A2(new_n294), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n212), .A2(new_n287), .ZN(new_n783));
  INV_X1    g0583(.A(new_n230), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n294), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(G20), .B1(KEYINPUT94), .B2(G169), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(KEYINPUT94), .A2(G169), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n252), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n776), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n209), .A2(new_n359), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n378), .A3(G200), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT95), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT95), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G303), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n378), .A2(new_n307), .A3(G190), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n359), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G326), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n806), .A2(new_n618), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n209), .A2(G190), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(new_n378), .A3(new_n307), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n811), .B1(G329), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n378), .A2(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n287), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n812), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(G311), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n812), .A2(new_n378), .A3(G200), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n807), .A2(G190), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n824), .A2(G283), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n803), .A2(new_n815), .A3(new_n822), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n823), .A2(new_n401), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n282), .B1(new_n820), .B2(new_n412), .C1(new_n222), .C2(new_n817), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(G50), .C2(new_n808), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n802), .A2(G87), .ZN(new_n832));
  INV_X1    g0632(.A(G159), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n813), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT32), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n831), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n805), .A2(G97), .B1(new_n825), .B2(G68), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT96), .Z(new_n838));
  OAI21_X1  g0638(.A(new_n828), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n796), .B1(new_n839), .B2(new_n790), .ZN(new_n840));
  INV_X1    g0640(.A(new_n793), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n708), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n778), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT97), .ZN(G396));
  OAI21_X1  g0644(.A(new_n418), .B1(new_n417), .B2(new_n706), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n415), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n415), .A2(new_n705), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n734), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n848), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n694), .A2(new_n706), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n768), .A2(G330), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n776), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n850), .A2(new_n792), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n790), .A2(new_n791), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n776), .B1(new_n859), .B2(G77), .ZN(new_n860));
  INV_X1    g0660(.A(new_n817), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G143), .A2(new_n861), .B1(new_n821), .B2(G159), .ZN(new_n862));
  INV_X1    g0662(.A(new_n825), .ZN(new_n863));
  INV_X1    g0663(.A(G150), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n862), .B1(new_n863), .B2(new_n864), .C1(new_n865), .C2(new_n809), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT34), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n282), .B1(new_n823), .B2(new_n325), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n806), .A2(new_n222), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n869), .B(new_n870), .C1(G132), .C2(new_n814), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n868), .B(new_n871), .C1(new_n202), .C2(new_n801), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n866), .A2(new_n867), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n809), .A2(new_n474), .B1(new_n820), .B2(new_n218), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G283), .B2(new_n825), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT99), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n823), .A2(new_n602), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n287), .B1(new_n817), .B2(new_n618), .C1(new_n806), .C2(new_n224), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n878), .B(new_n879), .C1(G311), .C2(new_n814), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n877), .B(new_n880), .C1(new_n401), .C2(new_n801), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n874), .B1(KEYINPUT100), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(KEYINPUT100), .B2(new_n881), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n857), .B(new_n860), .C1(new_n883), .C2(new_n790), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n856), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(G384));
  NOR2_X1   g0686(.A1(new_n773), .A2(new_n208), .ZN(new_n887));
  INV_X1    g0687(.A(G330), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n757), .A2(new_n762), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n756), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n760), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n451), .A2(new_n450), .A3(G169), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n445), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n434), .B(new_n705), .C1(new_n659), .C2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n453), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(KEYINPUT102), .A3(new_n434), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n434), .A2(new_n705), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n897), .A2(new_n457), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n848), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT103), .B1(new_n334), .B2(new_n338), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n342), .A2(new_n905), .A3(new_n343), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n906), .A3(new_n324), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n371), .B1(new_n907), .B2(new_n374), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n703), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n396), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n702), .B1(new_n380), .B2(new_n383), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n368), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n386), .A2(new_n389), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n386), .A2(new_n702), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n368), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT38), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n918), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(KEYINPUT104), .A3(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n902), .A2(new_n903), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n924), .ZN(new_n927));
  INV_X1    g0727(.A(new_n915), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n396), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT105), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT105), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n396), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n914), .A2(new_n915), .A3(new_n368), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n917), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n927), .B1(new_n936), .B2(new_n921), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n891), .A2(new_n901), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT40), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n926), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT107), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n459), .A2(new_n891), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT108), .Z(new_n943));
  AOI21_X1  g0743(.A(new_n888), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT106), .B1(new_n736), .B2(new_n459), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n734), .A2(new_n735), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n730), .A2(new_n731), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n684), .A2(new_n675), .A3(new_n558), .ZN(new_n949));
  AND4_X1   g0749(.A1(new_n505), .A2(new_n649), .A3(new_n510), .A4(new_n507), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n613), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(KEYINPUT29), .B(new_n706), .C1(new_n948), .C2(new_n951), .ZN(new_n952));
  AND4_X1   g0752(.A1(KEYINPUT106), .A2(new_n947), .A3(new_n459), .A4(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n665), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n851), .A2(new_n847), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n895), .A2(new_n900), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n955), .A2(new_n922), .A3(new_n925), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n658), .A2(new_n703), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n936), .A2(new_n921), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n924), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n897), .A2(new_n898), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n706), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n957), .B(new_n958), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n954), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n887), .B1(new_n945), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n945), .ZN(new_n969));
  INV_X1    g0769(.A(new_n528), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n218), .B(new_n232), .C1(new_n970), .C2(KEYINPUT35), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(KEYINPUT35), .B2(new_n970), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT36), .ZN(new_n973));
  OAI21_X1  g0773(.A(G77), .B1(new_n222), .B2(new_n325), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n230), .A2(new_n974), .B1(G50), .B2(new_n325), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n975), .A2(G1), .A3(new_n772), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT101), .Z(new_n978));
  NAND2_X1  g0778(.A1(new_n969), .A2(new_n978), .ZN(G367));
  OAI21_X1  g0779(.A(new_n571), .B1(new_n536), .B2(new_n706), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n689), .A2(new_n692), .A3(new_n705), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n714), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n705), .A2(new_n672), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n688), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n613), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n985), .B(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n983), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n684), .B1(new_n991), .B2(new_n649), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n706), .ZN(new_n993));
  INV_X1    g0793(.A(new_n982), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n716), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n993), .A2(new_n996), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n990), .B(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n720), .B(KEYINPUT41), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n718), .A2(new_n994), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n718), .A2(new_n994), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT111), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(new_n714), .ZN(new_n1009));
  MUX2_X1   g0809(.A(new_n713), .B(new_n711), .S(new_n715), .Z(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(new_n709), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n769), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1008), .A2(new_n714), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1009), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n999), .B1(new_n1015), .B2(new_n769), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n998), .B1(new_n1016), .B2(new_n775), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n242), .A2(new_n783), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n794), .B1(new_n212), .B2(new_n407), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n776), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n802), .A2(G58), .ZN(new_n1021));
  INV_X1    g0821(.A(G143), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n809), .A2(new_n1022), .B1(new_n823), .B2(new_n412), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G137), .B2(new_n814), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n282), .B1(new_n817), .B2(new_n864), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G50), .B2(new_n821), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n806), .A2(new_n325), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G159), .B2(new_n825), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1021), .A2(new_n1024), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n801), .A2(new_n218), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT46), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n287), .B1(new_n817), .B2(new_n474), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G283), .B2(new_n821), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n823), .A2(new_n224), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G311), .B2(new_n808), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n825), .A2(G294), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n814), .A2(G317), .B1(G107), .B2(new_n805), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT47), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1020), .B1(new_n1040), .B2(new_n790), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n841), .B2(new_n988), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1017), .A2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n713), .A2(new_n793), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n779), .A2(new_n721), .B1(G107), .B2(new_n212), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n239), .A2(new_n294), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n721), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n1047), .C1(G68), .C2(G77), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n405), .A2(new_n202), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT50), .Z(new_n1050));
  AOI21_X1  g0850(.A(new_n783), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1045), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n776), .B1(new_n1052), .B2(new_n795), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n282), .B1(new_n814), .B2(G326), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G317), .A2(new_n861), .B1(new_n821), .B2(G303), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n825), .A2(G311), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n818), .C2(new_n809), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT48), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n802), .A2(G294), .B1(G283), .B2(new_n805), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1054), .B1(new_n218), .B2(new_n823), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n861), .A2(G50), .B1(new_n408), .B2(new_n805), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT112), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n802), .A2(G77), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n287), .B(new_n1034), .C1(G68), .C2(new_n821), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n814), .A2(G150), .B1(G159), .B2(new_n808), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n347), .A2(new_n825), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1064), .A2(new_n1065), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1053), .B1(new_n1073), .B2(new_n790), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1011), .A2(new_n775), .B1(new_n1044), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1012), .A2(new_n771), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1011), .A2(new_n769), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(G393));
  NAND2_X1  g0881(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n774), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n249), .A2(new_n783), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n794), .B1(new_n224), .B2(new_n212), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n776), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n983), .A2(new_n841), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n813), .A2(new_n1022), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n806), .A2(new_n412), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G50), .C2(new_n825), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n287), .B(new_n878), .C1(new_n405), .C2(new_n821), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n325), .C2(new_n801), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n861), .A2(G159), .B1(G150), .B2(new_n808), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n861), .A2(G311), .B1(G317), .B2(new_n808), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n863), .A2(new_n474), .B1(new_n813), .B2(new_n818), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G116), .B2(new_n805), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n282), .B(new_n829), .C1(G294), .C2(new_n821), .ZN(new_n1099));
  INV_X1    g0899(.A(G283), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n801), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1092), .A2(new_n1094), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1086), .B(new_n1087), .C1(new_n790), .C2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1082), .A2(new_n1012), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n771), .A3(new_n1015), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(KEYINPUT118), .B1(new_n942), .B2(new_n888), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT118), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n459), .A2(new_n891), .A3(new_n1109), .A4(G330), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n665), .B(new_n1111), .C1(new_n946), .C2(new_n953), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n848), .A2(new_n888), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n891), .A2(new_n956), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n768), .A2(new_n1113), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n956), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n891), .A2(new_n1119), .A3(new_n956), .A4(new_n1113), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n768), .A2(new_n956), .A3(new_n1113), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n706), .B(new_n846), .C1(new_n948), .C2(new_n951), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n847), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n956), .B1(new_n891), .B2(new_n1113), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1121), .A2(new_n955), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n956), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT115), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT114), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n965), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n964), .A2(KEYINPUT114), .A3(new_n706), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n960), .A2(new_n924), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1117), .B1(new_n1123), .B2(new_n847), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n929), .A2(KEYINPUT105), .B1(new_n917), .B2(new_n934), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT38), .B1(new_n1138), .B2(new_n932), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1137), .B1(new_n1139), .B2(new_n927), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT115), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n955), .A2(new_n956), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n965), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n963), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1142), .B(new_n1145), .C1(new_n1147), .C2(new_n1122), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1130), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1136), .A2(new_n1140), .A3(KEYINPUT115), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT116), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1128), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n720), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1128), .A2(new_n1154), .A3(new_n1148), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1148), .A3(new_n775), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n776), .B1(new_n859), .B2(new_n347), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n863), .A2(new_n401), .B1(new_n813), .B2(new_n618), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G283), .B2(new_n808), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n287), .B1(new_n820), .B2(new_n224), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G116), .B2(new_n861), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1089), .B1(G68), .B2(new_n824), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n832), .A2(new_n1162), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n802), .A2(G150), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT53), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n863), .A2(new_n865), .B1(new_n823), .B2(new_n202), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G125), .B2(new_n814), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n282), .B1(new_n820), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G132), .B2(new_n861), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n805), .A2(G159), .B1(new_n808), .B2(G128), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1170), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1166), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1160), .B1(new_n1176), .B2(new_n790), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n963), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n792), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1158), .A2(new_n1159), .A3(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT120), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n311), .A2(new_n703), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n322), .B2(new_n421), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n421), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1186), .B(new_n1183), .C1(new_n313), .C2(new_n321), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1185), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n312), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n319), .B1(new_n318), .B2(new_n320), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n421), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1183), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n322), .A2(new_n421), .A3(new_n1184), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n940), .B2(G330), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n888), .B(new_n1197), .C1(new_n926), .C2(new_n939), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n966), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n957), .A2(new_n958), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n965), .B1(new_n959), .B2(new_n962), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n925), .A2(new_n903), .A3(new_n922), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n891), .B(new_n901), .C1(new_n1139), .C2(new_n927), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n902), .A2(new_n1205), .B1(new_n1206), .B2(KEYINPUT40), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1197), .B1(new_n1207), .B2(new_n888), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n940), .A2(G330), .A3(new_n1198), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1204), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1182), .B1(new_n1201), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n966), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1208), .A2(new_n1204), .A3(new_n1209), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(KEYINPUT120), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1112), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1211), .A2(new_n1214), .B1(new_n1215), .B2(new_n1157), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1181), .B1(new_n1216), .B2(KEYINPUT57), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1157), .A2(new_n1215), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1212), .A2(KEYINPUT120), .A3(new_n1213), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT120), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(KEYINPUT121), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1201), .A2(new_n1210), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(new_n1222), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n720), .B1(new_n1225), .B2(new_n1218), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1217), .A2(new_n1223), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1197), .A2(new_n791), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n282), .A2(G41), .ZN(new_n1229));
  AOI211_X1 g1029(.A(G50), .B(new_n1229), .C1(new_n327), .C2(new_n293), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1229), .B1(new_n407), .B2(new_n820), .C1(new_n401), .C2(new_n817), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1027), .B(new_n1231), .C1(G283), .C2(new_n814), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n823), .A2(new_n222), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n809), .A2(new_n218), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(G97), .C2(new_n825), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1068), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT58), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1230), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G128), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n817), .A2(new_n1239), .B1(new_n820), .B2(new_n865), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G132), .B2(new_n825), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n805), .A2(G150), .B1(new_n808), .B2(G125), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n801), .C2(new_n1171), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n327), .B(new_n293), .C1(new_n823), .C2(new_n833), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G124), .B2(new_n814), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1238), .B1(new_n1237), .B2(new_n1236), .C1(new_n1244), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n790), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT119), .Z(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n858), .A2(new_n202), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1228), .A2(new_n776), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1255), .B1(new_n1256), .B2(new_n775), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1227), .A2(new_n1257), .ZN(G375));
  OAI21_X1  g1058(.A(new_n776), .B1(new_n859), .B2(G68), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n808), .A2(G132), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n817), .B2(new_n865), .C1(new_n863), .C2(new_n1171), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n287), .B(new_n1233), .C1(G150), .C2(new_n821), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n814), .A2(G128), .B1(G50), .B2(new_n805), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n833), .C2(new_n801), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1264), .B2(KEYINPUT122), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(KEYINPUT122), .B2(new_n1264), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n802), .A2(G97), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n809), .A2(new_n618), .B1(new_n813), .B2(new_n474), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G116), .B2(new_n825), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n287), .B1(new_n820), .B2(new_n401), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G283), .B2(new_n861), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n824), .A2(G77), .B1(new_n408), .B2(new_n805), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1267), .A2(new_n1269), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1266), .A2(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(KEYINPUT123), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n790), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n1274), .B2(KEYINPUT123), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1259), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n956), .B2(new_n792), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1127), .B2(new_n774), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1280), .B(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1128), .A2(new_n999), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1112), .A2(new_n1127), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(G381));
  INV_X1    g1086(.A(G396), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1079), .A2(new_n1287), .A3(new_n1080), .ZN(new_n1288));
  OR4_X1    g1088(.A1(G384), .A2(G390), .A3(new_n1288), .A4(G381), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G387), .A2(new_n1289), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n704), .A2(G213), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G407), .B(G213), .C1(G375), .C2(new_n1294), .ZN(G409));
  NAND3_X1  g1095(.A1(new_n1227), .A2(G378), .A3(new_n1257), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1254), .B1(new_n774), .B2(new_n1224), .C1(new_n1221), .C2(new_n999), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1292), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1284), .B1(new_n1128), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1112), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n771), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1282), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n885), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1282), .A3(G384), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(KEYINPUT126), .A3(new_n1307), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1293), .A2(G2897), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1307), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1304), .B2(new_n1282), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1311), .B(new_n1309), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1300), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(G387), .A2(new_n1106), .A3(new_n1104), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(G390), .A2(new_n1017), .A3(new_n1042), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1288), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1287), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1319), .A2(new_n1324), .A3(new_n1320), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1329), .B1(new_n1300), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1293), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1333), .A2(KEYINPUT63), .A3(new_n1330), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1318), .A2(new_n1328), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1333), .A2(new_n1336), .A3(new_n1330), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1333), .B2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1336), .B1(new_n1333), .B2(new_n1330), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1337), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1335), .B1(new_n1342), .B2(new_n1328), .ZN(G405));
  NAND2_X1  g1143(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1291), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1296), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1348), .A2(new_n1330), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1326), .A2(new_n1327), .A3(KEYINPUT127), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1331), .B1(new_n1347), .B2(new_n1296), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1346), .A2(new_n1351), .A3(new_n1352), .A4(new_n1354), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1344), .B(new_n1345), .C1(new_n1350), .C2(new_n1353), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(G402));
endmodule


