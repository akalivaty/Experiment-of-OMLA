

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n420), .B(n302), .ZN(n303) );
  INV_X1 U320 ( .A(KEYINPUT87), .ZN(n400) );
  NOR2_X1 U321 ( .A1(n518), .A2(n461), .ZN(n566) );
  XOR2_X1 U322 ( .A(n307), .B(n306), .Z(n479) );
  XNOR2_X1 U323 ( .A(n396), .B(KEYINPUT28), .ZN(n535) );
  XOR2_X1 U324 ( .A(n385), .B(n384), .Z(n287) );
  XOR2_X1 U325 ( .A(n381), .B(G204GAT), .Z(n288) );
  XOR2_X1 U326 ( .A(KEYINPUT82), .B(KEYINPUT22), .Z(n289) );
  XOR2_X1 U327 ( .A(n452), .B(n451), .Z(n290) );
  XOR2_X1 U328 ( .A(G43GAT), .B(G50GAT), .Z(n291) );
  XOR2_X1 U329 ( .A(n433), .B(n379), .Z(n292) );
  XNOR2_X1 U330 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U331 ( .A(n301), .B(G85GAT), .ZN(n302) );
  XNOR2_X1 U332 ( .A(n429), .B(n428), .ZN(n431) );
  INV_X1 U333 ( .A(KEYINPUT54), .ZN(n459) );
  XNOR2_X1 U334 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U335 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U336 ( .A(n437), .B(n436), .ZN(n438) );
  NOR2_X1 U337 ( .A1(n516), .A2(n484), .ZN(n441) );
  NOR2_X1 U338 ( .A1(n465), .A2(n532), .ZN(n467) );
  XNOR2_X1 U339 ( .A(n467), .B(n466), .ZN(n561) );
  XOR2_X1 U340 ( .A(KEYINPUT94), .B(n442), .Z(n499) );
  XNOR2_X1 U341 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U342 ( .A(n443), .B(G29GAT), .ZN(n444) );
  XNOR2_X1 U343 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n445), .B(n444), .ZN(G1328GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n294) );
  XNOR2_X1 U346 ( .A(KEYINPUT74), .B(KEYINPUT9), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT10), .B(G92GAT), .Z(n296) );
  XNOR2_X1 U349 ( .A(G162GAT), .B(G106GAT), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n307) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n299), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U354 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n291), .B(n300), .ZN(n420) );
  AND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XOR2_X1 U357 ( .A(n348), .B(n303), .Z(n305) );
  XOR2_X1 U358 ( .A(G29GAT), .B(G134GAT), .Z(n321) );
  XOR2_X1 U359 ( .A(G99GAT), .B(KEYINPUT70), .Z(n434) );
  XNOR2_X1 U360 ( .A(n321), .B(n434), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U362 ( .A(KEYINPUT36), .B(n479), .ZN(n579) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U364 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n309) );
  NAND2_X1 U365 ( .A1(G231GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U367 ( .A(G8GAT), .B(G183GAT), .Z(n339) );
  XOR2_X1 U368 ( .A(n310), .B(n339), .Z(n318) );
  XOR2_X1 U369 ( .A(G78GAT), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U370 ( .A(G127GAT), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U372 ( .A(KEYINPUT12), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U373 ( .A(G1GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U375 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n417), .B(n319), .ZN(n320) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n427) );
  XOR2_X1 U379 ( .A(n320), .B(n427), .Z(n556) );
  INV_X1 U380 ( .A(n556), .ZN(n575) );
  XOR2_X1 U381 ( .A(KEYINPUT0), .B(G127GAT), .Z(n360) );
  XOR2_X1 U382 ( .A(n321), .B(n360), .Z(n323) );
  NAND2_X1 U383 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U385 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n325) );
  XNOR2_X1 U386 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U388 ( .A(n327), .B(n326), .Z(n333) );
  XOR2_X1 U389 ( .A(G113GAT), .B(G1GAT), .Z(n419) );
  XOR2_X1 U390 ( .A(KEYINPUT3), .B(G162GAT), .Z(n329) );
  XNOR2_X1 U391 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U393 ( .A(G141GAT), .B(n330), .Z(n386) );
  INV_X1 U394 ( .A(n386), .ZN(n331) );
  XOR2_X1 U395 ( .A(n419), .B(n331), .Z(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U397 ( .A(n334), .B(KEYINPUT1), .Z(n338) );
  XOR2_X1 U398 ( .A(G57GAT), .B(G85GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G120GAT), .B(G148GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n432) );
  XNOR2_X1 U401 ( .A(n432), .B(KEYINPUT5), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n397) );
  XOR2_X1 U403 ( .A(KEYINPUT86), .B(n339), .Z(n341) );
  NAND2_X1 U404 ( .A1(G226GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n356) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(G204GAT), .ZN(n347) );
  INV_X1 U407 ( .A(G92GAT), .ZN(n342) );
  NAND2_X1 U408 ( .A1(n342), .A2(G64GAT), .ZN(n345) );
  INV_X1 U409 ( .A(G64GAT), .ZN(n343) );
  NAND2_X1 U410 ( .A1(n343), .A2(G92GAT), .ZN(n344) );
  NAND2_X1 U411 ( .A1(n345), .A2(n344), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n425) );
  XOR2_X1 U413 ( .A(n348), .B(n425), .Z(n354) );
  XOR2_X1 U414 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n350) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n364) );
  XOR2_X1 U417 ( .A(G211GAT), .B(KEYINPUT80), .Z(n352) );
  XNOR2_X1 U418 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n382) );
  XNOR2_X1 U420 ( .A(n364), .B(n382), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n521) );
  XOR2_X1 U423 ( .A(G134GAT), .B(G190GAT), .Z(n358) );
  XNOR2_X1 U424 ( .A(G43GAT), .B(G99GAT), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U426 ( .A(n360), .B(n359), .Z(n362) );
  NAND2_X1 U427 ( .A1(G227GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U429 ( .A(n363), .B(G71GAT), .Z(n366) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(n364), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U432 ( .A(G120GAT), .B(G176GAT), .Z(n368) );
  XNOR2_X1 U433 ( .A(G113GAT), .B(G183GAT), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U435 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n370) );
  XNOR2_X1 U436 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U438 ( .A(n372), .B(n371), .Z(n373) );
  XOR2_X1 U439 ( .A(n374), .B(n373), .Z(n390) );
  AND2_X1 U440 ( .A1(n521), .A2(n390), .ZN(n375) );
  XOR2_X1 U441 ( .A(KEYINPUT88), .B(n375), .Z(n387) );
  XOR2_X1 U442 ( .A(KEYINPUT24), .B(G148GAT), .Z(n377) );
  XNOR2_X1 U443 ( .A(G22GAT), .B(KEYINPUT81), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U445 ( .A(G106GAT), .B(G78GAT), .Z(n433) );
  XNOR2_X1 U446 ( .A(G50GAT), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n289), .B(n378), .ZN(n379) );
  NAND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n292), .B(n380), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(KEYINPUT23), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n288), .B(n383), .ZN(n384) );
  XOR2_X1 U452 ( .A(n386), .B(n287), .Z(n462) );
  NAND2_X1 U453 ( .A1(n387), .A2(n462), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n388), .B(KEYINPUT25), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n389), .B(KEYINPUT89), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n521), .B(KEYINPUT27), .ZN(n398) );
  INV_X1 U457 ( .A(n390), .ZN(n532) );
  INV_X1 U458 ( .A(n532), .ZN(n524) );
  NOR2_X1 U459 ( .A1(n462), .A2(n524), .ZN(n391) );
  XOR2_X1 U460 ( .A(n391), .B(KEYINPUT26), .Z(n549) );
  INV_X1 U461 ( .A(n549), .ZN(n565) );
  NAND2_X1 U462 ( .A1(n398), .A2(n565), .ZN(n392) );
  NAND2_X1 U463 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U464 ( .A1(n397), .A2(n394), .ZN(n395) );
  XNOR2_X1 U465 ( .A(KEYINPUT90), .B(n395), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n462), .B(KEYINPUT65), .ZN(n396) );
  XNOR2_X1 U467 ( .A(KEYINPUT85), .B(n397), .ZN(n518) );
  NAND2_X1 U468 ( .A1(n398), .A2(n518), .ZN(n529) );
  NOR2_X1 U469 ( .A1(n535), .A2(n529), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n399), .A2(n532), .ZN(n401) );
  NAND2_X1 U471 ( .A1(n403), .A2(n402), .ZN(n482) );
  NAND2_X1 U472 ( .A1(n575), .A2(n482), .ZN(n404) );
  NOR2_X1 U473 ( .A1(n579), .A2(n404), .ZN(n405) );
  XNOR2_X1 U474 ( .A(KEYINPUT37), .B(n405), .ZN(n516) );
  XOR2_X1 U475 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n407) );
  NAND2_X1 U476 ( .A1(G229GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U477 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U478 ( .A(n408), .B(KEYINPUT66), .Z(n416) );
  XOR2_X1 U479 ( .A(G141GAT), .B(G29GAT), .Z(n410) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G36GAT), .ZN(n409) );
  XNOR2_X1 U481 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n412) );
  XNOR2_X1 U483 ( .A(G197GAT), .B(G8GAT), .ZN(n411) );
  XNOR2_X1 U484 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U485 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n418) );
  XOR2_X1 U487 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U488 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U489 ( .A(n422), .B(n421), .Z(n567) );
  INV_X1 U490 ( .A(n567), .ZN(n562) );
  XOR2_X1 U491 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n424) );
  XNOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT73), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n439) );
  XOR2_X1 U494 ( .A(n425), .B(KEYINPUT31), .Z(n429) );
  NAND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U496 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n437) );
  XOR2_X1 U498 ( .A(n433), .B(n432), .Z(n435) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n571) );
  NAND2_X1 U500 ( .A1(n562), .A2(n571), .ZN(n484) );
  XNOR2_X1 U501 ( .A(KEYINPUT95), .B(KEYINPUT38), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U503 ( .A1(n499), .A2(n518), .ZN(n445) );
  XOR2_X1 U504 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n443) );
  XNOR2_X1 U505 ( .A(n571), .B(KEYINPUT41), .ZN(n470) );
  NAND2_X1 U506 ( .A1(n470), .A2(n562), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n446), .B(KEYINPUT46), .ZN(n448) );
  INV_X1 U508 ( .A(n479), .ZN(n558) );
  NOR2_X1 U509 ( .A1(n558), .A2(n556), .ZN(n447) );
  AND2_X1 U510 ( .A1(n448), .A2(n447), .ZN(n450) );
  XNOR2_X1 U511 ( .A(KEYINPUT108), .B(KEYINPUT47), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n452) );
  NOR2_X1 U514 ( .A1(n575), .A2(n579), .ZN(n451) );
  NAND2_X1 U515 ( .A1(n571), .A2(n290), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n453), .B(KEYINPUT109), .ZN(n454) );
  NAND2_X1 U517 ( .A1(n454), .A2(n567), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n456), .A2(n455), .ZN(n457) );
  XOR2_X1 U519 ( .A(KEYINPUT48), .B(n457), .Z(n530) );
  XNOR2_X1 U520 ( .A(KEYINPUT117), .B(n521), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n530), .A2(n458), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U523 ( .A1(n566), .A2(n462), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U526 ( .A(KEYINPUT119), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n561), .A2(n556), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(G1350GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT99), .B(n470), .Z(n538) );
  NAND2_X1 U531 ( .A1(n561), .A2(n538), .ZN(n474) );
  XOR2_X1 U532 ( .A(G176GAT), .B(KEYINPUT57), .Z(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(G1349GAT) );
  NAND2_X1 U536 ( .A1(n561), .A2(n558), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n476) );
  XNOR2_X1 U538 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n475) );
  XOR2_X1 U539 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT76), .B(KEYINPUT16), .Z(n481) );
  NAND2_X1 U541 ( .A1(n556), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n483) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n501) );
  NOR2_X1 U544 ( .A1(n484), .A2(n501), .ZN(n493) );
  NAND2_X1 U545 ( .A1(n493), .A2(n518), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n521), .A2(n493), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT35), .B(KEYINPUT93), .Z(n490) );
  NAND2_X1 U551 ( .A1(n493), .A2(n524), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n492) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT92), .Z(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n493), .A2(n535), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT97), .Z(n496) );
  NAND2_X1 U558 ( .A1(n499), .A2(n521), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n524), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U563 ( .A1(n499), .A2(n535), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n567), .A2(n538), .ZN(n515) );
  NOR2_X1 U566 ( .A1(n501), .A2(n515), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(KEYINPUT100), .ZN(n511) );
  NAND2_X1 U568 ( .A1(n511), .A2(n518), .ZN(n506) );
  XOR2_X1 U569 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n504) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(KEYINPUT98), .B(n507), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U575 ( .A1(n511), .A2(n521), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n511), .A2(n524), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n513) );
  NAND2_X1 U580 ( .A1(n535), .A2(n511), .ZN(n512) );
  XNOR2_X1 U581 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(n514), .ZN(G1335GAT) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U585 ( .A(KEYINPUT105), .B(n517), .Z(n526) );
  NAND2_X1 U586 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U588 ( .A(G92GAT), .B(KEYINPUT107), .Z(n523) );
  NAND2_X1 U589 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n526), .A2(n535), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT112), .ZN(n537) );
  NOR2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(KEYINPUT110), .B(n531), .Z(n550) );
  NOR2_X1 U599 ( .A1(n550), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT111), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n562), .A2(n546), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U605 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n541), .Z(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n545) );
  XOR2_X1 U609 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U610 ( .A1(n546), .A2(n556), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U614 ( .A1(n546), .A2(n558), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n552) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n562), .A2(n559), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U621 ( .A1(n559), .A2(n470), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n556), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n578) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n578), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n578), .ZN(n576) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(n576), .Z(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(n580), .Z(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

