//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G141gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G148gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n203), .A2(new_n205), .B1(KEYINPUT2), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT79), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT80), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(G155gat), .B2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n206), .A2(KEYINPUT80), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(KEYINPUT80), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G155gat), .B2(G162gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(G155gat), .A3(G162gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n207), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n206), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(new_n208), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n226));
  NAND2_X1  g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(KEYINPUT22), .ZN(new_n229));
  INV_X1    g028(.A(G204gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G197gat), .ZN(new_n232));
  INV_X1    g031(.A(G197gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT74), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(KEYINPUT74), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(G197gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(G204gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n229), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G211gat), .A2(G218gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n227), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT75), .B1(new_n228), .B2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n226), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n228), .A2(KEYINPUT22), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n236), .A2(new_n237), .A3(G204gat), .ZN(new_n248));
  AOI21_X1  g047(.A(G204gat), .B1(new_n236), .B2(new_n237), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n243), .A2(new_n244), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT76), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n241), .A2(new_n227), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT77), .A3(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n254), .B(new_n247), .C1(new_n248), .C2(new_n249), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n225), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n246), .A2(new_n252), .B1(new_n255), .B2(new_n258), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n263), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n224), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G228gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n219), .B2(new_n223), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT82), .ZN(new_n271));
  INV_X1    g070(.A(new_n207), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n216), .B1(new_n214), .B2(new_n217), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n222), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n269), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT29), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n253), .A2(new_n259), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n268), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n276), .B2(new_n269), .ZN(new_n285));
  INV_X1    g084(.A(new_n269), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT82), .B(new_n286), .C1(new_n275), .C2(new_n222), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n263), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n235), .A2(new_n238), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n254), .B1(new_n290), .B2(new_n247), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n255), .B2(new_n258), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n269), .B1(new_n292), .B2(KEYINPUT29), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n219), .B2(new_n223), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n275), .A2(KEYINPUT83), .A3(new_n222), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  AOI211_X1 g097(.A(KEYINPUT86), .B(new_n268), .C1(new_n289), .C2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n300));
  INV_X1    g099(.A(new_n291), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT77), .B1(new_n239), .B2(new_n254), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n256), .A2(new_n257), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n286), .B1(new_n304), .B2(new_n284), .ZN(new_n305));
  INV_X1    g104(.A(new_n297), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n305), .A2(new_n306), .B1(new_n279), .B2(new_n280), .ZN(new_n307));
  INV_X1    g106(.A(new_n268), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n300), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n283), .B1(new_n299), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G22gat), .ZN(new_n311));
  INV_X1    g110(.A(G22gat), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n283), .B(new_n312), .C1(new_n299), .C2(new_n309), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT31), .B(G50gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT85), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT87), .B1(new_n263), .B2(KEYINPUT29), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n280), .A2(new_n261), .A3(new_n284), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(new_n225), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n281), .B1(new_n324), .B2(new_n224), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n288), .A2(new_n263), .B1(new_n293), .B2(new_n297), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(new_n326), .B2(new_n268), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n300), .A3(new_n308), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT89), .A3(new_n312), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT88), .B1(new_n329), .B2(new_n312), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n310), .A2(new_n333), .A3(G22gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n317), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n319), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n317), .B1(new_n311), .B2(KEYINPUT88), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n330), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n334), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT90), .A3(new_n319), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n344));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G134gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G127gat), .ZN(new_n349));
  INV_X1    g148(.A(G127gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G134gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(G113gat), .B2(G120gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G113gat), .A2(G120gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n352), .A2(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n351), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT72), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n345), .A2(KEYINPUT72), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT71), .B(G113gat), .Z(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n364), .B2(G120gat), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n347), .A2(new_n358), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n366), .B1(KEYINPUT3), .B2(new_n224), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n285), .B2(new_n287), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n276), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n295), .A2(new_n366), .A3(new_n296), .A4(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n347), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n363), .A2(new_n365), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n225), .B2(new_n276), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n271), .B2(new_n278), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n295), .A2(new_n366), .A3(new_n296), .A4(KEYINPUT4), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n371), .B1(new_n379), .B2(new_n224), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n375), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n224), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n369), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(KEYINPUT84), .A3(new_n224), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT5), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n376), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n376), .C1(new_n386), .C2(new_n392), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n368), .A2(new_n375), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT5), .B(new_n391), .C1(new_n403), .C2(new_n384), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n397), .B1(new_n404), .B2(new_n376), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(KEYINPUT23), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT66), .B(G176gat), .Z(new_n410));
  INV_X1    g209(.A(G169gat), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n411), .A2(KEYINPUT23), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G183gat), .A2(G190gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT24), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT65), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n413), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n427));
  NAND2_X1  g226(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n414), .A2(new_n425), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n417), .B(new_n418), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n411), .A2(KEYINPUT23), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT25), .B1(new_n432), .B2(G176gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(new_n409), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n423), .A2(new_n424), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n407), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT26), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n408), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n407), .A2(KEYINPUT26), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n414), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(KEYINPUT27), .B(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(KEYINPUT28), .A3(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n440), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n284), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g249(.A(G226gat), .B(G233gat), .C1(new_n435), .C2(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n263), .ZN(new_n453));
  XNOR2_X1  g252(.A(G8gat), .B(G36gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(G64gat), .B(G92gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n451), .A3(new_n280), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT30), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(KEYINPUT30), .A3(new_n456), .A4(new_n457), .ZN(new_n461));
  INV_X1    g260(.A(new_n456), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n450), .A2(new_n451), .A3(new_n280), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n280), .B1(new_n450), .B2(new_n451), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n406), .A2(new_n460), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n339), .A2(new_n343), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  INV_X1    g271(.A(new_n447), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n423), .A2(new_n424), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n431), .A2(new_n434), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n379), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n366), .B1(new_n435), .B2(new_n447), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G227gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n267), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n472), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT34), .B(new_n480), .C1(new_n476), .C2(new_n477), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT33), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G15gat), .B(G43gat), .Z(new_n489));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n485), .B(KEYINPUT32), .C1(new_n487), .C2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n484), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n482), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n492), .A2(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n492), .A2(new_n494), .ZN(new_n501));
  INV_X1    g300(.A(new_n484), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT73), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n492), .A3(new_n494), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n504), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n500), .B1(new_n507), .B2(KEYINPUT36), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT37), .B1(new_n463), .B2(new_n464), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n453), .A2(new_n510), .A3(new_n457), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n462), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n458), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT92), .B(new_n397), .C1(new_n404), .C2(new_n376), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n393), .B2(new_n398), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n400), .A2(new_n401), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n520), .A2(new_n521), .B1(KEYINPUT6), .B2(new_n405), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n460), .A2(new_n465), .A3(new_n461), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n393), .A2(new_n398), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT92), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n393), .A2(new_n518), .A3(new_n398), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n375), .B1(new_n368), .B2(new_n373), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n398), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n528), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n389), .A2(new_n390), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n529), .B1(new_n532), .B2(new_n375), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT40), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n539), .B(new_n530), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n516), .A2(new_n522), .B1(new_n527), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n508), .B1(new_n542), .B2(new_n337), .ZN(new_n543));
  INV_X1    g342(.A(new_n470), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n337), .A2(new_n544), .A3(new_n507), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n499), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n521), .A3(new_n526), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n523), .B1(new_n549), .B2(new_n399), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n550), .B2(KEYINPUT93), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n522), .B2(new_n523), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n553), .A3(new_n337), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n471), .A2(new_n543), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(KEYINPUT95), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT96), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n556), .B(new_n560), .ZN(new_n561));
  OAI22_X1  g360(.A1(new_n559), .A2(G1gat), .B1(KEYINPUT16), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n559), .A2(G1gat), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n562), .A2(new_n563), .A3(G8gat), .ZN(new_n564));
  OAI21_X1  g363(.A(G8gat), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G36gat), .ZN(new_n567));
  AND2_X1   g366(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(KEYINPUT17), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n565), .A3(new_n564), .ZN(new_n582));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n583), .B(KEYINPUT13), .Z(new_n587));
  NOR2_X1   g386(.A1(new_n566), .A2(new_n579), .ZN(new_n588));
  INV_X1    g387(.A(new_n579), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n564), .B2(new_n565), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT18), .A4(new_n583), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G197gat), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT11), .B(G169gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT94), .B(KEYINPUT12), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n599), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n586), .A2(new_n591), .A3(new_n601), .A4(new_n592), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n555), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT97), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n612));
  AND2_X1   g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G127gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n610), .B(KEYINPUT98), .Z(new_n616));
  AOI21_X1  g415(.A(new_n566), .B1(KEYINPUT21), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G155gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT7), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G99gat), .B(G106gat), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n631), .A2(new_n635), .A3(new_n633), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n637), .A2(KEYINPUT100), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(KEYINPUT100), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n581), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT101), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n645));
  AND2_X1   g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(KEYINPUT41), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n642), .B(new_n647), .C1(new_n589), .C2(new_n641), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n646), .A2(KEYINPUT41), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n653), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n610), .B1(new_n639), .B2(new_n640), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n638), .B1(new_n637), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n634), .B2(new_n636), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n611), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n616), .A2(KEYINPUT10), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n641), .ZN(new_n665));
  INV_X1    g464(.A(G230gat), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n663), .A2(new_n665), .B1(new_n666), .B2(new_n267), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n658), .A2(new_n662), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n267), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g470(.A(G120gat), .B(G148gat), .Z(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT105), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n673), .B(new_n674), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n670), .A3(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n626), .A2(new_n656), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n605), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n406), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(G1gat), .Z(G1324gat));
  NAND3_X1  g482(.A1(new_n605), .A2(new_n523), .A3(new_n680), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n684), .A2(G8gat), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT106), .B(KEYINPUT16), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G8gat), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(KEYINPUT42), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g489(.A(new_n508), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n681), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n499), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n681), .B2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n339), .A2(new_n343), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n656), .ZN(new_n700));
  INV_X1    g499(.A(new_n679), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n626), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n604), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n555), .A2(new_n700), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n406), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n571), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n555), .B2(new_n700), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n471), .A2(new_n543), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT73), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n499), .B2(new_n504), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n470), .B(new_n712), .C1(new_n342), .C2(new_n319), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n554), .B1(new_n713), .B2(new_n547), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n656), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n704), .B1(new_n709), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n406), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n708), .A2(new_n720), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n567), .A3(new_n523), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  INV_X1    g522(.A(new_n523), .ZN(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1329gat));
  AOI21_X1  g525(.A(G43gat), .B1(new_n705), .B2(new_n499), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n508), .A2(G43gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n718), .B2(new_n728), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(new_n337), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n718), .B2(new_n733), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n696), .A2(new_n702), .A3(G50gat), .A4(new_n700), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n605), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT48), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n337), .B(new_n704), .C1(new_n709), .C2(new_n717), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n732), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n696), .B(new_n704), .C1(new_n709), .C2(new_n717), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n736), .B1(new_n744), .B2(new_n732), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT109), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n736), .ZN(new_n748));
  INV_X1    g547(.A(new_n696), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n715), .B2(new_n656), .ZN(new_n751));
  INV_X1    g550(.A(new_n716), .ZN(new_n752));
  AOI211_X1 g551(.A(new_n700), .B(new_n752), .C1(new_n710), .C2(new_n714), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n749), .B(new_n703), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n748), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT48), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n743), .B1(new_n747), .B2(new_n757), .ZN(G1331gat));
  NOR4_X1   g557(.A1(new_n626), .A2(new_n656), .A3(new_n603), .A4(new_n701), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n715), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n406), .B(KEYINPUT111), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n760), .A2(new_n724), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  NOR3_X1   g568(.A1(new_n760), .A2(G71gat), .A3(new_n693), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(new_n508), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(G71gat), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n761), .A2(new_n749), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n625), .A2(new_n603), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n715), .A2(new_n656), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(new_n628), .A3(new_n706), .A4(new_n679), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n679), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n709), .B2(new_n717), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n706), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n628), .B2(new_n785), .ZN(G1336gat));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n523), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G92gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n777), .A2(new_n780), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n701), .A2(G92gat), .A3(new_n724), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n789), .B(new_n790), .C1(new_n777), .C2(new_n778), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n788), .B2(new_n791), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(G1337gat));
  INV_X1    g594(.A(G99gat), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n796), .A3(new_n499), .A4(new_n679), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n784), .A2(new_n508), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(new_n796), .ZN(G1338gat));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n733), .A2(new_n800), .A3(new_n679), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n789), .B(new_n802), .C1(new_n777), .C2(new_n778), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n784), .B2(new_n749), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n807));
  AND2_X1   g606(.A1(new_n784), .A2(new_n733), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n803), .B(new_n807), .C1(new_n808), .C2(new_n800), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1339gat));
  OR2_X1    g609(.A1(new_n588), .A2(new_n590), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n583), .B1(new_n580), .B2(new_n582), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n811), .A2(new_n587), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n597), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n602), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n664), .A2(new_n641), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n669), .C1(new_n668), .C2(new_n657), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n821), .B1(new_n666), .B2(new_n267), .C1(new_n663), .C2(new_n665), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n676), .A4(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n678), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n819), .A2(new_n667), .A3(KEYINPUT54), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n676), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n656), .A2(new_n817), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n828), .A2(new_n603), .A3(new_n678), .A4(new_n823), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n679), .A3(new_n602), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n656), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n626), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n680), .A2(new_n604), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n762), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n733), .A2(new_n712), .A3(new_n523), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n839), .A2(new_n364), .A3(new_n604), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n831), .A2(new_n832), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n700), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n829), .ZN(new_n843));
  AOI22_X1  g642(.A1(new_n843), .A2(new_n626), .B1(new_n604), .B2(new_n680), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n749), .A3(new_n693), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n406), .A2(new_n523), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n603), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(G113gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n848), .B2(G113gat), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(G1340gat));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n846), .ZN(new_n853));
  INV_X1    g652(.A(G120gat), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n701), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n679), .A3(new_n838), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n847), .A2(G127gat), .A3(new_n625), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT117), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n350), .B1(new_n839), .B2(new_n626), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n858), .A2(KEYINPUT117), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(G1342gat));
  NAND4_X1  g662(.A1(new_n837), .A2(new_n348), .A3(new_n656), .A4(new_n838), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT56), .Z(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n853), .B2(new_n700), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(KEYINPUT118), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(G1343gat));
  OAI21_X1  g668(.A(KEYINPUT57), .B1(new_n844), .B2(new_n696), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n836), .A2(new_n871), .A3(new_n733), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n691), .A2(new_n846), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n870), .A2(new_n603), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT119), .B1(new_n875), .B2(G141gat), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n508), .A2(new_n337), .A3(new_n523), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n604), .A2(G141gat), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n762), .A2(new_n836), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n879), .B1(new_n875), .B2(G141gat), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n876), .A2(new_n880), .A3(KEYINPUT58), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  AOI221_X4 g681(.A(new_n879), .B1(KEYINPUT119), .B2(new_n882), .C1(new_n875), .C2(G141gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n883), .ZN(G1344gat));
  NAND2_X1  g683(.A1(new_n837), .A2(new_n877), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n204), .A3(new_n679), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT59), .B(new_n204), .C1(new_n888), .C2(new_n679), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT57), .B1(new_n844), .B2(new_n337), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n836), .A2(new_n871), .A3(new_n749), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n891), .A2(new_n679), .A3(new_n892), .A4(new_n874), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n887), .B1(new_n889), .B2(new_n894), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n885), .A2(new_n626), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT120), .ZN(new_n897));
  AOI21_X1  g696(.A(G155gat), .B1(new_n896), .B2(KEYINPUT120), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n625), .A2(G155gat), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n897), .A2(new_n898), .B1(new_n888), .B2(new_n899), .ZN(G1346gat));
  INV_X1    g699(.A(G162gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n901), .A3(new_n656), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n888), .A2(new_n656), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n901), .ZN(G1347gat));
  INV_X1    g703(.A(new_n762), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(KEYINPUT121), .A3(new_n523), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n762), .B2(new_n724), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n845), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G169gat), .B1(new_n910), .B2(new_n604), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n706), .A2(new_n724), .ZN(new_n912));
  AND4_X1   g711(.A1(new_n337), .A2(new_n836), .A3(new_n507), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n411), .A3(new_n603), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT122), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n913), .B2(new_n679), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n845), .A2(new_n909), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n701), .A2(new_n410), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(G1349gat));
  OAI21_X1  g719(.A(G183gat), .B1(new_n910), .B2(new_n626), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n913), .A2(new_n441), .A3(new_n625), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g723(.A(new_n442), .B1(new_n918), .B2(new_n656), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n913), .A2(new_n442), .A3(new_n656), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n926), .A2(new_n929), .A3(new_n930), .ZN(G1351gat));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n691), .A3(new_n908), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n891), .A2(new_n892), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n233), .A3(new_n604), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n508), .A2(new_n337), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n836), .A2(new_n936), .A3(new_n912), .ZN(new_n937));
  AOI21_X1  g736(.A(G197gat), .B1(new_n937), .B2(new_n603), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n701), .A2(G204gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n836), .A2(new_n936), .A3(new_n912), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n934), .B2(new_n701), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1353gat));
  INV_X1    g747(.A(G211gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n937), .A2(new_n949), .A3(new_n625), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n891), .A2(new_n892), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n909), .A2(new_n691), .A3(new_n625), .ZN(new_n952));
  OAI21_X1  g751(.A(G211gat), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n700), .B1(new_n934), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n959), .B1(new_n958), .B2(new_n934), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G218gat), .ZN(new_n961));
  INV_X1    g760(.A(G218gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n937), .A2(new_n962), .A3(new_n656), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1355gat));
endmodule


