

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770;

  NOR2_X1 U366 ( .A1(n724), .A2(n637), .ZN(n636) );
  XNOR2_X1 U367 ( .A(KEYINPUT41), .B(n632), .ZN(n724) );
  XNOR2_X1 U368 ( .A(n646), .B(KEYINPUT38), .ZN(n696) );
  XNOR2_X1 U369 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  NAND2_X1 U370 ( .A1(n409), .A2(n408), .ZN(n345) );
  INV_X1 U371 ( .A(G116), .ZN(n494) );
  NOR2_X2 U372 ( .A1(n586), .A2(n486), .ZN(n357) );
  XOR2_X2 U373 ( .A(n663), .B(KEYINPUT62), .Z(n365) );
  INV_X2 U374 ( .A(KEYINPUT0), .ZN(n455) );
  NOR2_X2 U375 ( .A1(n593), .A2(KEYINPUT44), .ZN(n591) );
  XOR2_X2 U376 ( .A(n509), .B(n508), .Z(n366) );
  NOR2_X2 U377 ( .A1(n376), .A2(n374), .ZN(n659) );
  XNOR2_X2 U378 ( .A(n345), .B(n406), .ZN(n536) );
  NOR2_X1 U379 ( .A1(n707), .A2(n708), .ZN(n706) );
  BUF_X1 U380 ( .A(G116), .Z(n346) );
  NOR2_X1 U381 ( .A1(n596), .A2(n723), .ZN(n435) );
  NOR2_X2 U382 ( .A1(n700), .A2(n698), .ZN(n632) );
  INV_X1 U383 ( .A(n395), .ZN(n412) );
  NOR2_X1 U384 ( .A1(n618), .A2(n389), .ZN(n359) );
  XNOR2_X1 U385 ( .A(n539), .B(n444), .ZN(n710) );
  XNOR2_X1 U386 ( .A(n500), .B(KEYINPUT16), .ZN(n429) );
  XNOR2_X1 U387 ( .A(G134), .B(n346), .ZN(n569) );
  INV_X1 U388 ( .A(G122), .ZN(n500) );
  INV_X1 U389 ( .A(G113), .ZN(n495) );
  INV_X2 U390 ( .A(G953), .ZN(n759) );
  NAND2_X2 U391 ( .A1(n347), .A2(n481), .ZN(n425) );
  AND2_X1 U392 ( .A1(n347), .A2(n759), .ZN(n750) );
  XNOR2_X2 U393 ( .A(n484), .B(n367), .ZN(n347) );
  AND2_X1 U394 ( .A1(n443), .A2(n462), .ZN(n348) );
  BUF_X1 U395 ( .A(n445), .Z(n349) );
  XNOR2_X1 U396 ( .A(n489), .B(n488), .ZN(n445) );
  BUF_X1 U397 ( .A(n392), .Z(n350) );
  BUF_X1 U398 ( .A(n536), .Z(n351) );
  INV_X1 U399 ( .A(n425), .ZN(n352) );
  AND2_X2 U400 ( .A1(n425), .A2(n424), .ZN(n692) );
  INV_X1 U401 ( .A(G469), .ZN(n483) );
  INV_X1 U402 ( .A(G472), .ZN(n444) );
  NOR2_X1 U403 ( .A1(n663), .A2(G902), .ZN(n539) );
  XNOR2_X1 U404 ( .A(n375), .B(n363), .ZN(n374) );
  NOR2_X1 U405 ( .A1(n707), .A2(n617), .ZN(n633) );
  XNOR2_X1 U406 ( .A(n521), .B(n474), .ZN(n757) );
  XNOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n474) );
  XNOR2_X1 U408 ( .A(n464), .B(n463), .ZN(n723) );
  NAND2_X1 U409 ( .A1(n658), .A2(n389), .ZN(n388) );
  NOR2_X1 U410 ( .A1(n769), .A2(n770), .ZN(n375) );
  NOR2_X1 U411 ( .A1(G953), .A2(G237), .ZN(n550) );
  XNOR2_X1 U412 ( .A(n503), .B(n502), .ZN(n568) );
  XNOR2_X1 U413 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n502) );
  XNOR2_X1 U414 ( .A(n480), .B(G143), .ZN(n503) );
  INV_X1 U415 ( .A(G128), .ZN(n480) );
  XNOR2_X1 U416 ( .A(n568), .B(n504), .ZN(n510) );
  XNOR2_X1 U417 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n504) );
  OR2_X1 U418 ( .A1(G237), .A2(G902), .ZN(n542) );
  NAND2_X1 U419 ( .A1(n710), .A2(n695), .ZN(n380) );
  XOR2_X1 U420 ( .A(G101), .B(G146), .Z(n534) );
  XNOR2_X1 U421 ( .A(G131), .B(KEYINPUT5), .ZN(n533) );
  XNOR2_X1 U422 ( .A(n510), .B(n511), .ZN(n538) );
  XNOR2_X1 U423 ( .A(G137), .B(G134), .ZN(n511) );
  AND2_X1 U424 ( .A1(n469), .A2(n467), .ZN(n481) );
  INV_X1 U425 ( .A(n690), .ZN(n468) );
  XOR2_X1 U426 ( .A(G107), .B(G122), .Z(n570) );
  XNOR2_X1 U427 ( .A(n567), .B(n438), .ZN(n437) );
  INV_X1 U428 ( .A(KEYINPUT9), .ZN(n438) );
  XNOR2_X1 U429 ( .A(KEYINPUT101), .B(KEYINPUT99), .ZN(n439) );
  XNOR2_X1 U430 ( .A(KEYINPUT7), .B(KEYINPUT100), .ZN(n565) );
  XNOR2_X1 U431 ( .A(KEYINPUT88), .B(KEYINPUT72), .ZN(n466) );
  XNOR2_X1 U432 ( .A(n427), .B(n426), .ZN(n446) );
  XNOR2_X1 U433 ( .A(G101), .B(G110), .ZN(n426) );
  NAND2_X1 U434 ( .A1(n498), .A2(n499), .ZN(n427) );
  XNOR2_X1 U435 ( .A(n538), .B(n482), .ZN(n758) );
  XNOR2_X1 U436 ( .A(n557), .B(KEYINPUT87), .ZN(n482) );
  XNOR2_X1 U437 ( .A(n720), .B(n386), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n721), .B(KEYINPUT52), .ZN(n386) );
  INV_X1 U439 ( .A(n722), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n629), .B(KEYINPUT39), .ZN(n382) );
  NOR2_X1 U441 ( .A1(n682), .A2(n618), .ZN(n619) );
  XNOR2_X1 U442 ( .A(n575), .B(n440), .ZN(n595) );
  XNOR2_X1 U443 ( .A(KEYINPUT102), .B(G478), .ZN(n440) );
  NOR2_X1 U444 ( .A1(G902), .A2(n740), .ZN(n575) );
  INV_X1 U445 ( .A(KEYINPUT86), .ZN(n454) );
  XNOR2_X1 U446 ( .A(n529), .B(n530), .ZN(n743) );
  XNOR2_X1 U447 ( .A(n522), .B(n757), .ZN(n530) );
  XNOR2_X1 U448 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U449 ( .A1(n600), .A2(n708), .ZN(n487) );
  XNOR2_X1 U450 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n492) );
  XNOR2_X1 U451 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n493) );
  NAND2_X1 U452 ( .A1(n387), .A2(n712), .ZN(n713) );
  XNOR2_X1 U453 ( .A(n388), .B(KEYINPUT50), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n475), .B(G125), .ZN(n521) );
  INV_X1 U455 ( .A(G146), .ZN(n475) );
  XOR2_X1 U456 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n552) );
  XNOR2_X1 U457 ( .A(G143), .B(G113), .ZN(n558) );
  XNOR2_X1 U458 ( .A(G122), .B(G104), .ZN(n553) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n554) );
  INV_X1 U460 ( .A(n660), .ZN(n461) );
  XOR2_X1 U461 ( .A(G131), .B(G140), .Z(n557) );
  NAND2_X1 U462 ( .A1(n540), .A2(n660), .ZN(n541) );
  XNOR2_X1 U463 ( .A(G110), .B(G119), .ZN(n516) );
  XNOR2_X1 U464 ( .A(n526), .B(n525), .ZN(n528) );
  XNOR2_X1 U465 ( .A(G128), .B(G137), .ZN(n525) );
  NOR2_X1 U466 ( .A1(n419), .A2(n746), .ZN(n418) );
  NOR2_X1 U467 ( .A1(n432), .A2(G475), .ZN(n419) );
  INV_X1 U468 ( .A(KEYINPUT2), .ZN(n424) );
  INV_X1 U469 ( .A(KEYINPUT28), .ZN(n473) );
  AND2_X1 U470 ( .A1(n633), .A2(n710), .ZN(n634) );
  NOR2_X1 U471 ( .A1(n628), .A2(n627), .ZN(n644) );
  XNOR2_X1 U472 ( .A(n380), .B(n379), .ZN(n378) );
  INV_X1 U473 ( .A(KEYINPUT30), .ZN(n379) );
  XNOR2_X1 U474 ( .A(n538), .B(n372), .ZN(n663) );
  XNOR2_X1 U475 ( .A(n373), .B(n535), .ZN(n372) );
  XNOR2_X1 U476 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U477 ( .A(n761), .ZN(n371) );
  XNOR2_X1 U478 ( .A(n574), .B(n573), .ZN(n740) );
  XNOR2_X1 U479 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U480 ( .A(n437), .B(n354), .ZN(n574) );
  XNOR2_X1 U481 ( .A(n758), .B(n514), .ZN(n731) );
  XNOR2_X1 U482 ( .A(n512), .B(n466), .ZN(n465) );
  AND2_X1 U483 ( .A1(n383), .A2(n356), .ZN(n726) );
  NAND2_X1 U484 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U485 ( .A1(n382), .A2(n674), .ZN(n690) );
  AND2_X1 U486 ( .A1(n382), .A2(n381), .ZN(n631) );
  INV_X1 U487 ( .A(n630), .ZN(n381) );
  NOR2_X1 U488 ( .A1(n658), .A2(n657), .ZN(n688) );
  XNOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT35), .ZN(n589) );
  INV_X1 U490 ( .A(KEYINPUT32), .ZN(n488) );
  XNOR2_X1 U491 ( .A(n355), .B(n602), .ZN(n685) );
  OR2_X1 U492 ( .A1(n472), .A2(n470), .ZN(n680) );
  NAND2_X1 U493 ( .A1(n548), .A2(n635), .ZN(n470) );
  XNOR2_X1 U494 ( .A(n630), .B(KEYINPUT104), .ZN(n682) );
  XNOR2_X1 U495 ( .A(n532), .B(KEYINPUT25), .ZN(n476) );
  OR2_X1 U496 ( .A1(n743), .A2(G902), .ZN(n477) );
  AND2_X1 U497 ( .A1(n417), .A2(n416), .ZN(n415) );
  INV_X1 U498 ( .A(KEYINPUT56), .ZN(n433) );
  AND2_X1 U499 ( .A1(n418), .A2(KEYINPUT60), .ZN(n353) );
  XOR2_X1 U500 ( .A(n565), .B(n439), .Z(n354) );
  NOR2_X1 U501 ( .A1(n714), .A2(n453), .ZN(n355) );
  INV_X1 U502 ( .A(n521), .ZN(n448) );
  XOR2_X1 U503 ( .A(n725), .B(KEYINPUT116), .Z(n356) );
  AND2_X1 U504 ( .A1(G210), .A2(n542), .ZN(n358) );
  AND2_X1 U505 ( .A1(n420), .A2(n353), .ZN(n360) );
  NOR2_X1 U506 ( .A1(n705), .A2(n487), .ZN(n361) );
  XNOR2_X1 U507 ( .A(KEYINPUT34), .B(KEYINPUT74), .ZN(n362) );
  XOR2_X1 U508 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n363) );
  XNOR2_X1 U509 ( .A(KEYINPUT59), .B(KEYINPUT121), .ZN(n364) );
  INV_X1 U510 ( .A(n739), .ZN(n432) );
  XNOR2_X1 U511 ( .A(n738), .B(n364), .ZN(n739) );
  XNOR2_X1 U512 ( .A(KEYINPUT45), .B(KEYINPUT80), .ZN(n367) );
  AND2_X1 U513 ( .A1(n410), .A2(n430), .ZN(n368) );
  INV_X1 U514 ( .A(n422), .ZN(n421) );
  AND2_X1 U515 ( .A1(n739), .A2(n430), .ZN(n369) );
  NOR2_X1 U516 ( .A1(G952), .A2(n759), .ZN(n746) );
  INV_X1 U517 ( .A(n746), .ZN(n431) );
  INV_X1 U518 ( .A(KEYINPUT60), .ZN(n430) );
  NAND2_X1 U519 ( .A1(n590), .A2(n370), .ZN(n592) );
  XNOR2_X1 U520 ( .A(n370), .B(n767), .ZN(G24) );
  XNOR2_X2 U521 ( .A(n478), .B(n589), .ZN(n370) );
  XNOR2_X1 U522 ( .A(n481), .B(n371), .ZN(n760) );
  XNOR2_X1 U523 ( .A(n351), .B(n537), .ZN(n373) );
  NAND2_X1 U524 ( .A1(n377), .A2(n651), .ZN(n376) );
  INV_X1 U525 ( .A(n688), .ZN(n377) );
  NAND2_X1 U526 ( .A1(n378), .A2(n626), .ZN(n628) );
  NOR2_X1 U527 ( .A1(n731), .A2(G902), .ZN(n515) );
  INV_X1 U528 ( .A(n706), .ZN(n389) );
  BUF_X1 U529 ( .A(n501), .Z(n390) );
  OR2_X1 U530 ( .A1(n708), .A2(n610), .ZN(n391) );
  XNOR2_X2 U531 ( .A(n549), .B(n455), .ZN(n392) );
  XNOR2_X1 U532 ( .A(n549), .B(n455), .ZN(n582) );
  NAND2_X2 U533 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U534 ( .A1(n412), .A2(n418), .ZN(n411) );
  NAND2_X1 U535 ( .A1(n392), .A2(n581), .ZN(n393) );
  XNOR2_X1 U536 ( .A(n393), .B(n583), .ZN(n394) );
  XNOR2_X1 U537 ( .A(n584), .B(n583), .ZN(n402) );
  XNOR2_X1 U538 ( .A(n741), .B(n742), .ZN(n403) );
  XNOR2_X1 U539 ( .A(n735), .B(n736), .ZN(n404) );
  XNOR2_X1 U540 ( .A(n744), .B(n745), .ZN(n405) );
  NOR2_X2 U541 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X2 U542 ( .A1(n348), .A2(n456), .ZN(n395) );
  NAND2_X1 U543 ( .A1(n460), .A2(n456), .ZN(n737) );
  NAND2_X1 U544 ( .A1(n395), .A2(n421), .ZN(n420) );
  INV_X1 U545 ( .A(n692), .ZN(n459) );
  NAND2_X2 U546 ( .A1(n457), .A2(n459), .ZN(n456) );
  NAND2_X1 U547 ( .A1(n352), .A2(n398), .ZN(n396) );
  AND2_X2 U548 ( .A1(n396), .A2(n397), .ZN(n443) );
  OR2_X1 U549 ( .A1(KEYINPUT66), .A2(n461), .ZN(n397) );
  AND2_X1 U550 ( .A1(KEYINPUT2), .A2(n661), .ZN(n398) );
  INV_X1 U551 ( .A(n635), .ZN(n471) );
  BUF_X1 U552 ( .A(n653), .Z(n399) );
  BUF_X1 U553 ( .A(n401), .Z(n400) );
  NAND2_X1 U554 ( .A1(n423), .A2(KEYINPUT2), .ZN(n401) );
  NAND2_X1 U555 ( .A1(n357), .A2(n402), .ZN(n489) );
  NAND2_X1 U556 ( .A1(n394), .A2(n618), .ZN(n608) );
  AND2_X1 U557 ( .A1(n394), .A2(n361), .ZN(n673) );
  NOR2_X1 U558 ( .A1(n403), .A2(n746), .ZN(G63) );
  NOR2_X1 U559 ( .A1(n404), .A2(n746), .ZN(G54) );
  NOR2_X1 U560 ( .A1(n405), .A2(n746), .ZN(G66) );
  XNOR2_X2 U561 ( .A(G119), .B(KEYINPUT3), .ZN(n406) );
  NAND2_X1 U562 ( .A1(n495), .A2(G116), .ZN(n408) );
  NAND2_X1 U563 ( .A1(n494), .A2(G113), .ZN(n409) );
  XNOR2_X2 U564 ( .A(n536), .B(n429), .ZN(n428) );
  AND2_X2 U565 ( .A1(n401), .A2(n458), .ZN(n457) );
  NAND2_X1 U566 ( .A1(n693), .A2(n400), .ZN(n694) );
  NAND2_X1 U567 ( .A1(n411), .A2(n368), .ZN(n417) );
  NAND2_X1 U568 ( .A1(n422), .A2(n418), .ZN(n410) );
  NAND2_X1 U569 ( .A1(n360), .A2(n413), .ZN(n414) );
  NAND2_X1 U570 ( .A1(n412), .A2(n739), .ZN(n413) );
  NAND2_X1 U571 ( .A1(n415), .A2(n414), .ZN(G60) );
  NAND2_X1 U572 ( .A1(n412), .A2(n369), .ZN(n416) );
  NAND2_X1 U573 ( .A1(n432), .A2(G475), .ZN(n422) );
  INV_X1 U574 ( .A(n425), .ZN(n423) );
  XNOR2_X2 U575 ( .A(n428), .B(n446), .ZN(n501) );
  INV_X1 U576 ( .A(KEYINPUT66), .ZN(n661) );
  XNOR2_X1 U577 ( .A(n434), .B(n433), .ZN(G51) );
  NAND2_X1 U578 ( .A1(n436), .A2(n431), .ZN(n434) );
  XNOR2_X1 U579 ( .A(n435), .B(n362), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n662), .B(n366), .ZN(n436) );
  XNOR2_X2 U581 ( .A(n636), .B(KEYINPUT42), .ZN(n769) );
  NAND2_X1 U582 ( .A1(n441), .A2(n431), .ZN(n665) );
  XNOR2_X1 U583 ( .A(n664), .B(n365), .ZN(n441) );
  NAND2_X1 U584 ( .A1(n442), .A2(n603), .ZN(n604) );
  NAND2_X1 U585 ( .A1(n685), .A2(n668), .ZN(n442) );
  AND2_X1 U586 ( .A1(n606), .A2(n391), .ZN(n485) );
  NAND2_X1 U587 ( .A1(n705), .A2(n706), .ZN(n599) );
  AND2_X2 U588 ( .A1(n443), .A2(n462), .ZN(n460) );
  NOR2_X2 U589 ( .A1(n445), .A2(n673), .ZN(n587) );
  XNOR2_X1 U590 ( .A(n349), .B(n768), .ZN(G21) );
  XNOR2_X1 U591 ( .A(n446), .B(n465), .ZN(n513) );
  NAND2_X1 U592 ( .A1(n491), .A2(n490), .ZN(n451) );
  NAND2_X1 U593 ( .A1(n447), .A2(n491), .ZN(n452) );
  NOR2_X1 U594 ( .A1(n449), .A2(n448), .ZN(n447) );
  INV_X1 U595 ( .A(n490), .ZN(n449) );
  NAND2_X1 U596 ( .A1(n452), .A2(n450), .ZN(n507) );
  NAND2_X1 U597 ( .A1(n451), .A2(n448), .ZN(n450) );
  INV_X1 U598 ( .A(n350), .ZN(n453) );
  XNOR2_X1 U599 ( .A(n392), .B(n454), .ZN(n596) );
  NOR2_X1 U600 ( .A1(n660), .A2(n661), .ZN(n458) );
  NAND2_X1 U601 ( .A1(n692), .A2(n661), .ZN(n462) );
  NAND2_X1 U602 ( .A1(n705), .A2(n359), .ZN(n464) );
  INV_X1 U603 ( .A(KEYINPUT33), .ZN(n463) );
  NOR2_X1 U604 ( .A1(n766), .A2(n468), .ZN(n467) );
  XNOR2_X1 U605 ( .A(n659), .B(KEYINPUT48), .ZN(n469) );
  XNOR2_X1 U606 ( .A(n634), .B(n473), .ZN(n472) );
  OR2_X1 U607 ( .A1(n472), .A2(n471), .ZN(n637) );
  INV_X1 U608 ( .A(n680), .ZN(n675) );
  XNOR2_X2 U609 ( .A(n477), .B(n476), .ZN(n708) );
  NAND2_X1 U610 ( .A1(n479), .A2(n643), .ZN(n478) );
  XNOR2_X2 U611 ( .A(n635), .B(KEYINPUT1), .ZN(n705) );
  XNOR2_X2 U612 ( .A(n515), .B(n483), .ZN(n635) );
  XNOR2_X2 U613 ( .A(n653), .B(KEYINPUT19), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n607), .A2(n485), .ZN(n484) );
  INV_X1 U615 ( .A(n618), .ZN(n486) );
  NAND2_X1 U616 ( .A1(n501), .A2(n492), .ZN(n490) );
  OR2_X2 U617 ( .A1(n501), .A2(n493), .ZN(n491) );
  INV_X1 U618 ( .A(KEYINPUT24), .ZN(n518) );
  INV_X1 U619 ( .A(n707), .ZN(n579) );
  XNOR2_X1 U620 ( .A(n518), .B(KEYINPUT89), .ZN(n519) );
  AND2_X1 U621 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U622 ( .A(KEYINPUT90), .ZN(n527) );
  XNOR2_X1 U623 ( .A(n513), .B(G146), .ZN(n514) );
  XNOR2_X1 U624 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n583) );
  XNOR2_X1 U625 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n509) );
  INV_X1 U626 ( .A(G107), .ZN(n496) );
  NAND2_X1 U627 ( .A1(n496), .A2(G104), .ZN(n499) );
  INV_X1 U628 ( .A(G104), .ZN(n497) );
  NAND2_X1 U629 ( .A1(n497), .A2(G107), .ZN(n498) );
  NAND2_X1 U630 ( .A1(G224), .A2(n759), .ZN(n505) );
  XNOR2_X1 U631 ( .A(n510), .B(n505), .ZN(n506) );
  XNOR2_X2 U632 ( .A(n507), .B(n506), .ZN(n540) );
  XNOR2_X1 U633 ( .A(n540), .B(KEYINPUT84), .ZN(n508) );
  NAND2_X1 U634 ( .A1(G227), .A2(n759), .ZN(n512) );
  INV_X1 U635 ( .A(n705), .ZN(n658) );
  XOR2_X1 U636 ( .A(KEYINPUT23), .B(G140), .Z(n517) );
  XNOR2_X1 U637 ( .A(n517), .B(n516), .ZN(n520) );
  XNOR2_X1 U638 ( .A(n520), .B(n519), .ZN(n522) );
  XOR2_X1 U639 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n524) );
  NAND2_X1 U640 ( .A1(G234), .A2(n759), .ZN(n523) );
  XNOR2_X1 U641 ( .A(n524), .B(n523), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n566), .A2(G221), .ZN(n526) );
  NAND2_X1 U643 ( .A1(G234), .A2(n660), .ZN(n531) );
  XNOR2_X1 U644 ( .A(KEYINPUT20), .B(n531), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n576), .A2(G217), .ZN(n532) );
  NAND2_X1 U646 ( .A1(n550), .A2(G210), .ZN(n537) );
  INV_X1 U647 ( .A(n710), .ZN(n600) );
  XNOR2_X2 U648 ( .A(n541), .B(n358), .ZN(n623) );
  NAND2_X1 U649 ( .A1(G214), .A2(n542), .ZN(n695) );
  NAND2_X2 U650 ( .A1(n623), .A2(n695), .ZN(n653) );
  NAND2_X1 U651 ( .A1(G234), .A2(G237), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n543), .B(KEYINPUT14), .ZN(n544) );
  NAND2_X1 U653 ( .A1(G952), .A2(n544), .ZN(n722) );
  NOR2_X1 U654 ( .A1(G953), .A2(n722), .ZN(n615) );
  NAND2_X1 U655 ( .A1(G902), .A2(n544), .ZN(n611) );
  INV_X1 U656 ( .A(G898), .ZN(n749) );
  NAND2_X1 U657 ( .A1(G953), .A2(n749), .ZN(n752) );
  NOR2_X1 U658 ( .A1(n611), .A2(n752), .ZN(n545) );
  NOR2_X1 U659 ( .A1(n615), .A2(n545), .ZN(n546) );
  XNOR2_X1 U660 ( .A(KEYINPUT85), .B(n546), .ZN(n547) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n563) );
  NAND2_X1 U662 ( .A1(G214), .A2(n550), .ZN(n551) );
  XNOR2_X1 U663 ( .A(n552), .B(n551), .ZN(n556) );
  XNOR2_X1 U664 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U665 ( .A(n556), .B(n555), .Z(n561) );
  XNOR2_X1 U666 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U667 ( .A(n757), .B(n559), .ZN(n560) );
  XNOR2_X1 U668 ( .A(n561), .B(n560), .ZN(n738) );
  NOR2_X1 U669 ( .A1(G902), .A2(n738), .ZN(n562) );
  XNOR2_X1 U670 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U671 ( .A(G475), .B(n564), .Z(n594) );
  INV_X1 U672 ( .A(n594), .ZN(n588) );
  NAND2_X1 U673 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U674 ( .A(n568), .B(KEYINPUT98), .ZN(n572) );
  XNOR2_X1 U675 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U676 ( .A1(n588), .A2(n595), .ZN(n698) );
  INV_X1 U677 ( .A(n698), .ZN(n580) );
  XOR2_X1 U678 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n578) );
  NAND2_X1 U679 ( .A1(G221), .A2(n576), .ZN(n577) );
  XNOR2_X1 U680 ( .A(n578), .B(n577), .ZN(n707) );
  NAND2_X1 U681 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U682 ( .A(n710), .B(KEYINPUT6), .ZN(n618) );
  AND2_X1 U683 ( .A1(n705), .A2(n708), .ZN(n585) );
  XNOR2_X1 U684 ( .A(n585), .B(KEYINPUT103), .ZN(n586) );
  XNOR2_X1 U685 ( .A(n587), .B(KEYINPUT82), .ZN(n590) );
  NOR2_X1 U686 ( .A1(n595), .A2(n588), .ZN(n643) );
  INV_X1 U687 ( .A(KEYINPUT70), .ZN(n593) );
  XNOR2_X1 U688 ( .A(n592), .B(n591), .ZN(n607) );
  NAND2_X1 U689 ( .A1(n593), .A2(KEYINPUT44), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n595), .A2(n594), .ZN(n630) );
  NOR2_X1 U691 ( .A1(n595), .A2(n594), .ZN(n674) );
  INV_X1 U692 ( .A(n674), .ZN(n684) );
  NAND2_X1 U693 ( .A1(n630), .A2(n684), .ZN(n699) );
  XNOR2_X1 U694 ( .A(n699), .B(KEYINPUT78), .ZN(n603) );
  NAND2_X1 U695 ( .A1(n635), .A2(n706), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n596), .A2(n627), .ZN(n597) );
  XNOR2_X1 U697 ( .A(n597), .B(KEYINPUT92), .ZN(n598) );
  NAND2_X1 U698 ( .A1(n598), .A2(n600), .ZN(n668) );
  NOR2_X1 U699 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U700 ( .A(KEYINPUT93), .B(n601), .ZN(n714) );
  XNOR2_X1 U701 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n602) );
  AND2_X1 U702 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U703 ( .A1(n705), .A2(n608), .ZN(n609) );
  XNOR2_X1 U704 ( .A(n609), .B(KEYINPUT81), .ZN(n610) );
  NOR2_X1 U705 ( .A1(n708), .A2(n610), .ZN(n666) );
  NOR2_X1 U706 ( .A1(G900), .A2(n611), .ZN(n612) );
  NAND2_X1 U707 ( .A1(G953), .A2(n612), .ZN(n613) );
  XNOR2_X1 U708 ( .A(KEYINPUT105), .B(n613), .ZN(n614) );
  NOR2_X1 U709 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U710 ( .A(KEYINPUT76), .B(n616), .Z(n626) );
  NAND2_X1 U711 ( .A1(n626), .A2(n708), .ZN(n617) );
  NAND2_X1 U712 ( .A1(n633), .A2(n619), .ZN(n620) );
  XNOR2_X1 U713 ( .A(KEYINPUT106), .B(n620), .ZN(n654) );
  NOR2_X1 U714 ( .A1(n654), .A2(n705), .ZN(n621) );
  NAND2_X1 U715 ( .A1(n621), .A2(n695), .ZN(n622) );
  XNOR2_X1 U716 ( .A(n622), .B(KEYINPUT43), .ZN(n624) );
  INV_X1 U717 ( .A(n623), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n624), .A2(n646), .ZN(n625) );
  XNOR2_X1 U719 ( .A(KEYINPUT107), .B(n625), .ZN(n766) );
  NAND2_X1 U720 ( .A1(n644), .A2(n696), .ZN(n629) );
  XNOR2_X1 U721 ( .A(n631), .B(KEYINPUT40), .ZN(n770) );
  NAND2_X1 U722 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U723 ( .A1(KEYINPUT78), .A2(n680), .ZN(n638) );
  NOR2_X1 U724 ( .A1(KEYINPUT47), .A2(n638), .ZN(n639) );
  NOR2_X1 U725 ( .A1(n699), .A2(n639), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n680), .B(KEYINPUT47), .ZN(n642) );
  NAND2_X1 U727 ( .A1(KEYINPUT78), .A2(n699), .ZN(n640) );
  NAND2_X1 U728 ( .A1(n675), .A2(n640), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n678) );
  XNOR2_X1 U732 ( .A(KEYINPUT79), .B(n678), .ZN(n647) );
  NAND2_X1 U733 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U735 ( .A(KEYINPUT83), .B(KEYINPUT108), .ZN(n652) );
  XNOR2_X1 U736 ( .A(n652), .B(KEYINPUT36), .ZN(n656) );
  NOR2_X1 U737 ( .A1(n654), .A2(n399), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n737), .A2(G210), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n737), .A2(G472), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U742 ( .A(G101), .B(n666), .Z(G3) );
  NOR2_X1 U743 ( .A1(n682), .A2(n668), .ZN(n667) );
  XOR2_X1 U744 ( .A(G104), .B(n667), .Z(G6) );
  NOR2_X1 U745 ( .A1(n668), .A2(n684), .ZN(n672) );
  XOR2_X1 U746 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n670) );
  XNOR2_X1 U747 ( .A(G107), .B(KEYINPUT27), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U749 ( .A(n672), .B(n671), .ZN(G9) );
  XOR2_X1 U750 ( .A(G110), .B(n673), .Z(G12) );
  XOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .Z(n677) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n677), .B(n676), .ZN(G30) );
  XOR2_X1 U754 ( .A(G143), .B(n678), .Z(n679) );
  XNOR2_X1 U755 ( .A(KEYINPUT110), .B(n679), .ZN(G45) );
  NOR2_X1 U756 ( .A1(n682), .A2(n680), .ZN(n681) );
  XOR2_X1 U757 ( .A(G146), .B(n681), .Z(G48) );
  NOR2_X1 U758 ( .A1(n682), .A2(n685), .ZN(n683) );
  XOR2_X1 U759 ( .A(G113), .B(n683), .Z(G15) );
  NOR2_X1 U760 ( .A1(n685), .A2(n684), .ZN(n687) );
  XNOR2_X1 U761 ( .A(n346), .B(KEYINPUT111), .ZN(n686) );
  XNOR2_X1 U762 ( .A(n687), .B(n686), .ZN(G18) );
  XNOR2_X1 U763 ( .A(G125), .B(n688), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U765 ( .A(G134), .B(KEYINPUT112), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n691), .B(n690), .ZN(G36) );
  XNOR2_X1 U767 ( .A(n692), .B(KEYINPUT77), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n694), .A2(n759), .ZN(n728) );
  NOR2_X1 U769 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n703) );
  INV_X1 U771 ( .A(n699), .ZN(n701) );
  NOR2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U774 ( .A1(n723), .A2(n704), .ZN(n719) );
  NAND2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT49), .ZN(n711) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U779 ( .A(KEYINPUT51), .B(n715), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n724), .A2(n716), .ZN(n717) );
  XOR2_X1 U781 ( .A(KEYINPUT113), .B(n717), .Z(n718) );
  NOR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U783 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n721) );
  NOR2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U785 ( .A(n726), .B(KEYINPUT117), .ZN(n727) );
  XNOR2_X1 U786 ( .A(n729), .B(KEYINPUT118), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n730), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n733) );
  XNOR2_X1 U789 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n732) );
  XNOR2_X1 U790 ( .A(n733), .B(n732), .ZN(n734) );
  XOR2_X1 U791 ( .A(n731), .B(n734), .Z(n736) );
  NAND2_X1 U792 ( .A1(G469), .A2(n395), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n740), .B(KEYINPUT122), .ZN(n742) );
  NAND2_X1 U794 ( .A1(n395), .A2(G478), .ZN(n741) );
  XOR2_X1 U795 ( .A(n743), .B(KEYINPUT123), .Z(n745) );
  NAND2_X1 U796 ( .A1(G217), .A2(n395), .ZN(n744) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n747) );
  XOR2_X1 U798 ( .A(KEYINPUT61), .B(n747), .Z(n748) );
  NOR2_X1 U799 ( .A1(n749), .A2(n748), .ZN(n751) );
  NOR2_X1 U800 ( .A1(n751), .A2(n750), .ZN(n756) );
  XNOR2_X1 U801 ( .A(n390), .B(KEYINPUT124), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U803 ( .A(n754), .B(KEYINPUT125), .ZN(n755) );
  XOR2_X1 U804 ( .A(n756), .B(n755), .Z(G69) );
  XOR2_X1 U805 ( .A(n758), .B(n757), .Z(n761) );
  NAND2_X1 U806 ( .A1(n760), .A2(n759), .ZN(n765) );
  XNOR2_X1 U807 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n762), .A2(G900), .ZN(n763) );
  NAND2_X1 U809 ( .A1(n763), .A2(G953), .ZN(n764) );
  NAND2_X1 U810 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U811 ( .A(G140), .B(n766), .Z(G42) );
  XNOR2_X1 U812 ( .A(G122), .B(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U813 ( .A(G119), .B(KEYINPUT127), .ZN(n768) );
  XOR2_X1 U814 ( .A(n769), .B(G137), .Z(G39) );
  XOR2_X1 U815 ( .A(G131), .B(n770), .Z(G33) );
endmodule

