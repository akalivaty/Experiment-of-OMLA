//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n206));
  NAND4_X1  g005(.A1(new_n203), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT27), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n211), .A3(new_n204), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n206), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n217), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n207), .A2(new_n214), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT24), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(G169gat), .ZN(new_n225));
  INV_X1    g024(.A(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n204), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT24), .A3(new_n221), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n222), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n223), .ZN(new_n233));
  AND4_X1   g032(.A1(KEYINPUT25), .A2(new_n232), .A3(new_n233), .A4(new_n230), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n219), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(G113gat), .B2(G120gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n242), .B(KEYINPUT65), .C1(new_n238), .C2(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n244), .A2(new_n245), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(new_n219), .C1(new_n231), .C2(new_n234), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G227gat), .ZN(new_n251));
  INV_X1    g050(.A(G233gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT32), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n251), .A2(new_n252), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n247), .A2(new_n256), .A3(new_n249), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n247), .A2(new_n249), .A3(new_n259), .A4(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n255), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT33), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  XNOR2_X1  g061(.A(G15gat), .B(G43gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(G71gat), .B(G99gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n261), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT33), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n261), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n254), .B1(new_n266), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT34), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n258), .A2(new_n260), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n269), .ZN(new_n282));
  INV_X1    g081(.A(new_n265), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n254), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n272), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n274), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n279), .B1(new_n274), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n202), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n279), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n266), .A2(new_n273), .A3(new_n254), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n285), .B1(new_n284), .B2(new_n272), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n279), .A3(new_n286), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(KEYINPUT36), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296));
  INV_X1    g095(.A(G228gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n252), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n300));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301));
  XOR2_X1   g100(.A(G155gat), .B(G162gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n303), .A3(new_n306), .ZN(new_n308));
  XNOR2_X1  g107(.A(G155gat), .B(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  AND2_X1   g112(.A1(G211gat), .A2(G218gat), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(KEYINPUT22), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(G211gat), .A2(G218gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n315), .B(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n312), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n319), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n298), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n322), .B1(new_n320), .B2(KEYINPUT75), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n315), .B(new_n317), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n324), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n312), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n326), .A2(new_n298), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n327), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G22gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT3), .B1(new_n330), .B2(new_n331), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n331), .B2(new_n330), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n334), .B1(new_n340), .B2(new_n312), .ZN(new_n341));
  OAI21_X1  g140(.A(G22gat), .B1(new_n341), .B2(new_n327), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT74), .B(KEYINPUT31), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(G50gat), .ZN(new_n344));
  XOR2_X1   g143(.A(G78gat), .B(G106gat), .Z(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  AND4_X1   g145(.A1(new_n296), .A2(new_n338), .A3(new_n342), .A4(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT76), .B1(new_n336), .B2(new_n337), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n348), .A2(new_n346), .B1(new_n338), .B2(new_n342), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n355), .B(KEYINPUT70), .Z(new_n356));
  NAND2_X1  g155(.A1(new_n235), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n235), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT71), .B(new_n219), .C1(new_n231), .C2(new_n234), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n355), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n329), .B(new_n357), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n356), .B1(new_n235), .B2(new_n324), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n319), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n354), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n366), .A3(new_n354), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(KEYINPUT30), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n366), .ZN(new_n371));
  INV_X1    g170(.A(new_n354), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n371), .A2(KEYINPUT30), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n311), .A2(new_n246), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n304), .A2(new_n244), .A3(new_n310), .A4(new_n245), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n304), .A2(KEYINPUT3), .A3(new_n310), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n323), .A2(new_n248), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n377), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n311), .A2(new_n383), .A3(new_n246), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n311), .B2(new_n246), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT5), .B(new_n379), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n385), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n311), .A2(new_n383), .A3(new_n246), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n311), .A2(new_n246), .A3(KEYINPUT73), .A4(new_n383), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n378), .A2(KEYINPUT5), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n391), .A2(new_n381), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n396), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(G57gat), .B(G85gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n400), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n394), .A3(new_n399), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n370), .A2(new_n373), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n289), .A2(new_n295), .B1(new_n351), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n392), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n378), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n376), .A2(new_n378), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT39), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n413), .B(new_n378), .C1(new_n409), .C2(new_n410), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n399), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n415), .A2(KEYINPUT40), .A3(new_n399), .A4(new_n416), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n419), .A2(new_n402), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n373), .A4(new_n370), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT77), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n370), .A2(new_n373), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n402), .A3(new_n420), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n405), .A2(new_n401), .A3(new_n369), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT37), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n354), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n367), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n363), .B2(new_n366), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT38), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT38), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n319), .B(new_n357), .C1(new_n361), .C2(new_n362), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n329), .B1(new_n364), .B2(new_n365), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(KEYINPUT37), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n436), .C1(new_n367), .C2(new_n429), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n426), .A3(new_n438), .A4(new_n350), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n287), .A2(new_n288), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT35), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n350), .A4(new_n406), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n293), .A2(new_n350), .A3(new_n406), .A4(new_n294), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n408), .A2(new_n439), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT78), .B(G29gat), .ZN(new_n447));
  INV_X1    g246(.A(G36gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(G29gat), .A2(G36gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT14), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT15), .B(new_n446), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(KEYINPUT79), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n450), .B(KEYINPUT14), .Z(new_n457));
  OR2_X1    g256(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n452), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n464), .A2(G1gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n464), .B1(new_n466), .B2(G1gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(KEYINPUT80), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G8gat), .ZN(new_n469));
  INV_X1    g268(.A(G8gat), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT80), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT17), .B(new_n452), .C1(new_n456), .C2(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n463), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n471), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n461), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n476), .B2(new_n461), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n474), .B(new_n475), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n461), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT81), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n475), .A4(new_n474), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n482), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n482), .A2(KEYINPUT84), .A3(new_n488), .A4(new_n483), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(new_n475), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n480), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n476), .A2(new_n461), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n486), .A2(KEYINPUT18), .A3(new_n475), .A4(new_n474), .ZN(new_n498));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(G197gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT11), .B(G169gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT12), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n491), .A2(new_n492), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n497), .A3(new_n498), .ZN(new_n506));
  INV_X1    g305(.A(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n445), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G71gat), .B(G78gat), .Z(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT86), .ZN(new_n513));
  INV_X1    g312(.A(G57gat), .ZN(new_n514));
  INV_X1    g313(.A(G64gat), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT85), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n514), .B2(KEYINPUT85), .ZN(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n513), .A2(new_n518), .A3(new_n519), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G57gat), .B(G64gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n512), .B1(new_n524), .B2(new_n517), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT20), .ZN(new_n531));
  XNOR2_X1  g330(.A(G183gat), .B(G211gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n472), .B1(new_n527), .B2(new_n526), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT89), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT88), .ZN(new_n537));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n535), .B(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n540), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n546), .B2(new_n547), .ZN(new_n550));
  NAND3_X1  g349(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n544), .B1(new_n461), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(KEYINPUT90), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n461), .B2(new_n462), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n559), .A2(new_n560), .B1(new_n473), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n564), .ZN(new_n568));
  XNOR2_X1  g367(.A(G134gat), .B(G162gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n562), .B2(new_n564), .ZN(new_n573));
  INV_X1    g372(.A(new_n571), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n561), .A2(new_n473), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n563), .B(new_n575), .C1(new_n560), .C2(new_n559), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n573), .A2(new_n574), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n552), .B(new_n553), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT92), .B1(new_n583), .B2(new_n526), .ZN(new_n584));
  INV_X1    g383(.A(new_n556), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(new_n523), .A3(new_n554), .A4(new_n525), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT94), .ZN(new_n589));
  INV_X1    g388(.A(new_n526), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(KEYINPUT92), .A3(new_n557), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n582), .B1(new_n593), .B2(KEYINPUT95), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT10), .B1(new_n587), .B2(new_n591), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT10), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT93), .B1(new_n586), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n590), .A2(new_n599), .A3(new_n557), .A4(KEYINPUT10), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n595), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n594), .B(new_n602), .C1(KEYINPUT95), .C2(new_n593), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n592), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n582), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n543), .A2(new_n578), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n511), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n405), .A2(new_n401), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g412(.A1(new_n608), .A2(new_n424), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT96), .B(KEYINPUT16), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G8gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n470), .B2(new_n614), .ZN(new_n618));
  MUX2_X1   g417(.A(new_n617), .B(new_n618), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g418(.A1(new_n289), .A2(new_n295), .ZN(new_n620));
  OAI21_X1  g419(.A(G15gat), .B1(new_n608), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n440), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(G15gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n608), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT97), .ZN(G1326gat));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n350), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT98), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT43), .B(G22gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(G1327gat));
  NAND2_X1  g428(.A1(new_n541), .A2(new_n542), .ZN(new_n630));
  INV_X1    g429(.A(new_n578), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n630), .A2(new_n631), .A3(new_n606), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n511), .A2(new_n611), .A3(new_n447), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT45), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n445), .B2(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n442), .A2(new_n444), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n351), .A2(new_n407), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n287), .A2(new_n288), .A3(new_n202), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT36), .B1(new_n293), .B2(new_n294), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n439), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT44), .A3(new_n578), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n606), .B(KEYINPUT100), .Z(new_n648));
  NOR3_X1   g447(.A1(new_n648), .A2(new_n510), .A3(new_n630), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n610), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n636), .B(new_n637), .C1(new_n651), .C2(new_n447), .ZN(G1328gat));
  INV_X1    g451(.A(new_n424), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n647), .A2(new_n653), .A3(new_n649), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n448), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n511), .A2(new_n633), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n658), .A2(G36gat), .A3(new_n424), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT46), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(G1329gat));
  INV_X1    g460(.A(new_n620), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G43gat), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n658), .A2(new_n622), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n650), .A2(new_n663), .B1(G43gat), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g465(.A1(new_n639), .A2(new_n646), .A3(new_n351), .A4(new_n649), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT102), .B1(new_n667), .B2(G50gat), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT48), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n658), .A2(G50gat), .A3(new_n350), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(G50gat), .B2(new_n667), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n672), .ZN(G1331gat));
  INV_X1    g472(.A(new_n648), .ZN(new_n674));
  NOR4_X1   g473(.A1(new_n674), .A2(new_n543), .A3(new_n509), .A4(new_n578), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n645), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n645), .A2(KEYINPUT103), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n610), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(G57gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1332gat));
  AND2_X1   g482(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n424), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n688));
  OR2_X1    g487(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n687), .B2(new_n688), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(G1333gat));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n680), .B2(new_n622), .ZN(new_n694));
  INV_X1    g493(.A(G71gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n678), .A2(KEYINPUT106), .A3(new_n440), .A4(new_n679), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n684), .A2(G71gat), .A3(new_n662), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT50), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT50), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1334gat));
  NOR2_X1   g502(.A1(new_n680), .A2(new_n350), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT107), .B(G78gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1335gat));
  NOR2_X1   g505(.A1(new_n630), .A2(new_n509), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n606), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n647), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G85gat), .B1(new_n711), .B2(new_n610), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  NOR4_X1   g512(.A1(new_n445), .A2(new_n713), .A3(new_n631), .A4(new_n708), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n631), .B1(new_n640), .B2(new_n644), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT51), .B1(new_n715), .B2(new_n707), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n611), .A2(new_n546), .A3(new_n606), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n717), .B2(new_n718), .ZN(G1336gat));
  NOR3_X1   g518(.A1(new_n674), .A2(G92gat), .A3(new_n424), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n714), .B2(new_n716), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT109), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n639), .A2(new_n646), .A3(new_n653), .A4(new_n710), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT52), .B1(new_n723), .B2(G92gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n725), .B(new_n720), .C1(new_n714), .C2(new_n716), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n445), .A2(new_n631), .A3(new_n708), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n713), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n707), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n733), .A3(new_n720), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n723), .A2(G92gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n728), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT110), .B1(new_n727), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n724), .A3(new_n726), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n734), .A2(new_n735), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n728), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n711), .B2(new_n620), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n622), .A2(G99gat), .A3(new_n709), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n717), .B2(new_n744), .ZN(G1338gat));
  NOR3_X1   g544(.A1(new_n674), .A2(G106gat), .A3(new_n350), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n733), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT111), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n647), .A2(new_n351), .A3(new_n710), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G106gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n747), .A2(KEYINPUT111), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT53), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754));
  INV_X1    g553(.A(new_n746), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n750), .B(new_n754), .C1(new_n717), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(G1339gat));
  OR3_X1    g556(.A1(new_n596), .A2(new_n601), .A3(new_n595), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(KEYINPUT54), .A3(new_n602), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n760), .B(new_n595), .C1(new_n596), .C2(new_n601), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n582), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n761), .B2(new_n582), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(KEYINPUT55), .B(new_n759), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n509), .A2(new_n767), .A3(new_n603), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n494), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n486), .B(new_n770), .C1(new_n476), .C2(new_n461), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n475), .B1(new_n486), .B2(new_n474), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n502), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(KEYINPUT113), .B(new_n502), .C1(new_n772), .C2(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n505), .A3(new_n606), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n578), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n767), .A2(new_n578), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n505), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n768), .A2(new_n603), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n543), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n607), .A2(new_n510), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n351), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n653), .A2(new_n610), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n622), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n791), .A2(new_n236), .A3(new_n510), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n785), .A2(new_n786), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n622), .A2(new_n351), .ZN(new_n794));
  AND4_X1   g593(.A1(new_n611), .A2(new_n793), .A3(new_n424), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n509), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n236), .B2(new_n796), .ZN(G1340gat));
  OAI21_X1  g596(.A(G120gat), .B1(new_n791), .B2(new_n674), .ZN(new_n798));
  INV_X1    g597(.A(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n606), .A2(new_n237), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT114), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT115), .ZN(G1341gat));
  AOI21_X1  g602(.A(G127gat), .B1(new_n795), .B2(new_n630), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n787), .A2(G127gat), .A3(new_n630), .A4(new_n790), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(G1342gat));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n631), .A2(G134gat), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n795), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n810), .B1(new_n795), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT56), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n812), .A2(new_n813), .A3(KEYINPUT56), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n812), .C2(new_n813), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n791), .B2(new_n631), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n662), .A2(new_n789), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n793), .B2(new_n351), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n824), .B(new_n350), .C1(new_n785), .C2(new_n786), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n509), .B(new_n822), .C1(new_n823), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G141gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n620), .A2(new_n351), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n653), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n510), .A2(G141gat), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n793), .A2(new_n611), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n821), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n610), .B1(new_n785), .B2(new_n786), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(KEYINPUT119), .A3(new_n829), .A4(new_n830), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n821), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(G141gat), .B2(new_n826), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT120), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n837), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n827), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n829), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n826), .A2(G141gat), .B1(new_n844), .B2(new_n830), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n841), .B(new_n842), .C1(new_n821), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n839), .A2(new_n846), .ZN(G1344gat));
  OR3_X1    g646(.A1(new_n843), .A2(G148gat), .A3(new_n709), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n823), .A2(new_n825), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n606), .A3(new_n822), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(G148gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n851), .B2(G148gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(G1345gat));
  AOI21_X1  g654(.A(G155gat), .B1(new_n844), .B2(new_n630), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n849), .A2(new_n662), .A3(new_n789), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n630), .A2(G155gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT121), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(G1346gat));
  AOI21_X1  g659(.A(G162gat), .B1(new_n844), .B2(new_n578), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n578), .A2(G162gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(G1347gat));
  AOI21_X1  g662(.A(new_n611), .B1(new_n785), .B2(new_n786), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n864), .A2(new_n653), .A3(new_n794), .ZN(new_n865));
  AOI21_X1  g664(.A(G169gat), .B1(new_n865), .B2(new_n509), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n653), .A2(new_n610), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n622), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT122), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(new_n787), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n510), .A2(new_n225), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(G1348gat));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n226), .A3(new_n606), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n870), .A2(new_n648), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n226), .ZN(G1349gat));
  NAND3_X1  g674(.A1(new_n865), .A2(new_n203), .A3(new_n630), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n870), .A2(new_n630), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n208), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n865), .A2(new_n204), .A3(new_n578), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n870), .A2(new_n578), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G190gat), .ZN(new_n882));
  XOR2_X1   g681(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(G1351gat));
  NAND4_X1  g685(.A1(new_n620), .A2(KEYINPUT124), .A3(new_n653), .A4(new_n351), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n828), .B2(new_n424), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n864), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(G197gat), .B1(new_n890), .B2(new_n509), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n850), .A2(KEYINPUT125), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n849), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n662), .A2(new_n867), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n896), .A2(G197gat), .A3(new_n509), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n891), .B1(new_n895), .B2(new_n897), .ZN(G1352gat));
  XOR2_X1   g697(.A(KEYINPUT126), .B(G204gat), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n890), .A2(new_n606), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT62), .Z(new_n901));
  INV_X1    g700(.A(new_n896), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n674), .B(new_n902), .C1(new_n892), .C2(new_n894), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n903), .B2(new_n899), .ZN(G1353gat));
  INV_X1    g703(.A(G211gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n905), .A3(new_n630), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n896), .A2(new_n630), .ZN(new_n907));
  OAI21_X1  g706(.A(G211gat), .B1(new_n849), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  AOI21_X1  g711(.A(G218gat), .B1(new_n890), .B2(new_n578), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n578), .A2(G218gat), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT127), .Z(new_n915));
  NOR2_X1   g714(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n895), .B2(new_n916), .ZN(G1355gat));
endmodule


