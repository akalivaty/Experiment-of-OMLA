//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n445, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT68), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n463), .B2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(KEYINPUT70), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n460), .A2(new_n461), .ZN(new_n486));
  AND2_X1   g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(KEYINPUT71), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n460), .B2(new_n461), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n485), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n464), .A2(G138), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n486), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n464), .A2(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n462), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n492), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n506), .B1(new_n503), .B2(new_n504), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(G88), .B1(new_n507), .B2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n501), .A2(new_n502), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n509), .B2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(G89), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g101(.A(G51), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n521), .A2(new_n528), .ZN(G168));
  OAI211_X1 g104(.A(G52), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n515), .A2(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G64), .B1(new_n514), .B2(new_n515), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n509), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  XNOR2_X1  g112(.A(KEYINPUT6), .B(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G43), .A3(G543), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n531), .ZN(new_n541));
  OAI21_X1  g116(.A(G56), .B1(new_n514), .B2(new_n515), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n509), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(new_n507), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n507), .A2(new_n554), .A3(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n531), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n510), .A2(new_n538), .A3(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G91), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT74), .B(G65), .Z(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n516), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n556), .A2(new_n560), .A3(new_n564), .ZN(G299));
  OAI21_X1  g140(.A(KEYINPUT75), .B1(new_n533), .B2(new_n536), .ZN(new_n566));
  INV_X1    g141(.A(G64), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n501), .B2(new_n502), .ZN(new_n568));
  INV_X1    g143(.A(new_n535), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT72), .B(G90), .Z(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(new_n510), .A3(new_n538), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .A4(new_n530), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G301));
  INV_X1    g151(.A(G89), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n503), .B2(new_n504), .ZN(new_n578));
  INV_X1    g153(.A(new_n520), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n510), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n580), .A2(new_n527), .A3(new_n526), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n551), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n507), .A2(KEYINPUT76), .A3(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n558), .A2(G87), .A3(new_n559), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n558), .A2(G86), .A3(new_n559), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n516), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n507), .A2(G48), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n509), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n507), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n531), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n505), .A2(G85), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n602), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT78), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT80), .B(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n516), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n558), .A2(G92), .A3(new_n559), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(KEYINPUT79), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n558), .A2(new_n616), .A3(G92), .A4(new_n559), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n615), .B1(new_n614), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n608), .B1(G868), .B2(new_n621), .ZN(G284));
  OAI21_X1  g197(.A(new_n608), .B1(G868), .B2(new_n621), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n621), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n486), .A2(new_n465), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n463), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n477), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n464), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT81), .Z(G156));
  INV_X1    g222(.A(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT83), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n664), .A3(new_n666), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n665), .A2(new_n666), .ZN(new_n675));
  INV_X1    g250(.A(new_n664), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n668), .B1(new_n676), .B2(new_n667), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT84), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n684), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n692), .A2(new_n689), .A3(new_n684), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n690), .B1(new_n689), .B2(new_n684), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g280(.A1(G162), .A2(G29), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G29), .B2(G35), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(G2090), .ZN(new_n713));
  INV_X1    g288(.A(G2090), .ZN(new_n714));
  OAI211_X1 g289(.A(KEYINPUT99), .B(new_n714), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(new_n464), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n463), .A2(G139), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT25), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n717), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n723), .B2(G33), .ZN(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT93), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G20), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT101), .B(G1956), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n713), .A2(new_n715), .A3(new_n728), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n712), .A2(G2090), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G129), .B2(new_n477), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G32), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  NOR2_X1   g321(.A1(G164), .A2(new_n723), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G27), .B2(new_n723), .ZN(new_n748));
  INV_X1    g323(.A(G2078), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n723), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT96), .B1(new_n644), .B2(new_n723), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT97), .B(G28), .Z(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(KEYINPUT30), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT30), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(new_n723), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n753), .B(new_n754), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  NOR2_X1   g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n723), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT94), .Z(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n471), .B2(new_n723), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n725), .C2(new_n726), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n730), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n730), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n730), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n730), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G1966), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G1966), .ZN(new_n776));
  INV_X1    g351(.A(new_n771), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n769), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n737), .A2(new_n746), .A3(new_n760), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n736), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT89), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n620), .B2(new_n730), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT90), .B(G1348), .Z(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n730), .A2(G19), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n545), .B2(new_n730), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1341), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n723), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT91), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT28), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n463), .A2(G140), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n477), .A2(G128), .ZN(new_n796));
  OR2_X1    g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(new_n723), .ZN(new_n801));
  INV_X1    g376(.A(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n787), .A2(new_n788), .A3(new_n791), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n782), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT102), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n782), .A2(KEYINPUT102), .A3(new_n806), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT88), .Z(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n463), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n477), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(G29), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT87), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n816), .A2(new_n817), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n730), .A2(G22), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G166), .B2(new_n730), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1971), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n730), .A2(G23), .ZN(new_n832));
  AND3_X1   g407(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n730), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT33), .B(G1976), .Z(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G305), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n730), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G6), .B2(new_n730), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT32), .B(G1981), .Z(new_n841));
  AOI22_X1  g416(.A1(new_n840), .A2(new_n841), .B1(new_n834), .B2(new_n835), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n837), .B(new_n842), .C1(new_n840), .C2(new_n841), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n828), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n812), .A2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n812), .A2(new_n849), .ZN(G150));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n507), .A2(G55), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n510), .A2(new_n538), .A3(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(G67), .B1(new_n514), .B2(new_n515), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n509), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n853), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n860), .A2(KEYINPUT103), .A3(new_n509), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n852), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT103), .B1(new_n860), .B2(new_n509), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n853), .A2(new_n854), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n858), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT105), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n621), .A2(G559), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT106), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  INV_X1    g447(.A(new_n545), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n862), .A2(new_n873), .A3(new_n866), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n545), .B1(new_n859), .B2(new_n861), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n545), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n871), .B(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n875), .A2(new_n876), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT104), .B1(new_n878), .B2(new_n545), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G860), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n881), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n869), .B1(new_n891), .B2(new_n892), .ZN(G145));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n495), .A2(new_n894), .A3(new_n497), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n495), .B2(new_n497), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n492), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(new_n799), .ZN(new_n898));
  AOI22_X1  g473(.A1(G130), .A2(new_n477), .B1(new_n463), .B2(G142), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n900), .A2(new_n464), .A3(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n464), .B2(G118), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n902), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n898), .B(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n722), .B(new_n742), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n635), .B(new_n822), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n908), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n644), .B(new_n471), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(new_n481), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G37), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .A4(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n511), .A2(new_n509), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n507), .A2(G50), .ZN(new_n925));
  INV_X1    g500(.A(G88), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n531), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n923), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n508), .B(KEYINPUT110), .C1(new_n509), .C2(new_n511), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n833), .ZN(new_n931));
  NAND3_X1  g506(.A1(G288), .A2(new_n928), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(G290), .A2(new_n838), .ZN(new_n934));
  OAI211_X1 g509(.A(G305), .B(new_n598), .C1(new_n602), .C2(new_n605), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n931), .A2(new_n934), .A3(new_n935), .A4(new_n932), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n630), .B(new_n886), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n614), .A2(new_n617), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT10), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n625), .B1(new_n946), .B2(new_n612), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n625), .B(new_n612), .C1(new_n618), .C2(new_n619), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n947), .B2(new_n949), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n620), .A2(G299), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(KEYINPUT41), .A3(new_n948), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n942), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n941), .A2(new_n952), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n941), .B1(new_n952), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G868), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n867), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(G295));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n961), .A2(new_n965), .A3(new_n963), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n961), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(G331));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n969));
  NOR2_X1   g544(.A1(KEYINPUT43), .A2(G37), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n566), .A2(new_n574), .A3(G168), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(G171), .B2(G286), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n566), .A2(new_n574), .A3(new_n972), .A4(G168), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n886), .A2(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n566), .A2(G168), .A3(new_n574), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n570), .A2(new_n530), .A3(new_n573), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(new_n979), .B2(G168), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n880), .A2(new_n981), .A3(new_n874), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n954), .A2(new_n956), .A3(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n977), .A2(new_n955), .A3(new_n982), .A4(new_n948), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n939), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n970), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n954), .A2(new_n983), .A3(new_n956), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n939), .B1(new_n988), .B2(new_n985), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n969), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n914), .B1(new_n984), .B2(new_n986), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n991), .B2(new_n989), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n985), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n937), .A2(new_n938), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n970), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n880), .A2(new_n981), .A3(new_n874), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n981), .B1(new_n874), .B2(new_n880), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(new_n950), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n1000), .B2(new_n988), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n995), .A2(new_n1001), .A3(KEYINPUT113), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n990), .A2(new_n992), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n991), .B2(new_n989), .ZN(new_n1006));
  AOI21_X1  g581(.A(G37), .B1(new_n1000), .B2(new_n988), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n995), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(KEYINPUT43), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1004), .B1(new_n995), .B2(new_n1001), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1005), .A2(new_n1012), .A3(KEYINPUT115), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(G397));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(G1966), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n897), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n466), .A2(G40), .A3(new_n470), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(G1384), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1023), .B1(G164), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n499), .A2(new_n1020), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1022), .B1(new_n1031), .B2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n897), .A2(new_n1033), .A3(new_n1020), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n766), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT121), .B(new_n1019), .C1(new_n1021), .C2(new_n1027), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1030), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT118), .B(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G168), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1018), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1039), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT51), .B(new_n1040), .C1(new_n1037), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT124), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(new_n1045), .A3(new_n1040), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1045), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1042), .A2(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT62), .ZN(new_n1051));
  OAI221_X1 g626(.A(new_n1051), .B1(new_n1047), .B2(new_n1048), .C1(new_n1042), .C2(new_n1044), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G303), .A2(G8), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT55), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1022), .B1(new_n897), .B2(new_n1025), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1031), .A2(new_n1024), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1971), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1058), .A2(KEYINPUT117), .B1(new_n1059), .B2(G2090), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1058), .A2(KEYINPUT117), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1055), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n897), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1043), .C1(new_n1064), .C2(G288), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n590), .A2(new_n1069), .A3(new_n594), .A4(new_n595), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(KEYINPUT120), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(KEYINPUT120), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n505), .A2(G86), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n594), .A2(new_n595), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G1981), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT49), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1063), .A2(new_n1043), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(KEYINPUT49), .A3(new_n1076), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1065), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1079), .A2(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1023), .B1(new_n1031), .B2(KEYINPUT50), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1033), .B1(new_n897), .B2(new_n1020), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1058), .B1(new_n714), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1054), .B1(new_n1087), .B2(new_n1039), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1062), .A2(new_n1068), .A3(new_n1083), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1090), .B1(new_n1091), .B2(G2078), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1059), .A2(new_n778), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(G2078), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1092), .B(new_n1093), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n575), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1050), .A2(new_n1052), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1102));
  XOR2_X1   g677(.A(G299), .B(KEYINPUT57), .Z(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1056), .A2(new_n1057), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1348), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1063), .A2(G2067), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n620), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1103), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1111), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1106), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1106), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1111), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1109), .A2(KEYINPUT60), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1109), .A2(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n621), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1114), .B(new_n1117), .C1(new_n1118), .C2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT58), .B(G1341), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1063), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1091), .B2(G1996), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n545), .ZN(new_n1125));
  NAND2_X1  g700(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1127), .B(new_n1128), .C1(new_n621), .C2(new_n1119), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1112), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1022), .B(new_n1096), .C1(new_n897), .C2(new_n1025), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1021), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1092), .A2(new_n1093), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G301), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT54), .B1(new_n1135), .B2(new_n1098), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1089), .ZN(new_n1137));
  OAI221_X1 g712(.A(KEYINPUT54), .B1(new_n1097), .B2(new_n575), .C1(new_n979), .C2(new_n1134), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1130), .A2(new_n1137), .A3(new_n1049), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1068), .A2(new_n1083), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G288), .A2(G1976), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1140), .A2(new_n1062), .B1(new_n1143), .B2(new_n1078), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1068), .A2(new_n1083), .A3(KEYINPUT63), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1037), .A2(G168), .A3(new_n1043), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(G8), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1054), .A2(KEYINPUT122), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1145), .A2(new_n1147), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1089), .B2(new_n1146), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1144), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1100), .A2(new_n1139), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n822), .B(new_n826), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT116), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n799), .B(new_n802), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n742), .B(G1996), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(G290), .B(G1986), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1159), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1157), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1158), .A2(G1996), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT46), .Z(new_n1171));
  OAI21_X1  g746(.A(new_n1159), .B1(new_n742), .B2(new_n1163), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n822), .A2(new_n826), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1165), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n800), .A2(new_n802), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1158), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1158), .A2(G1986), .A3(G290), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT126), .Z(new_n1183));
  INV_X1    g758(.A(KEYINPUT48), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1183), .A2(new_n1184), .B1(new_n1159), .B2(new_n1166), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1181), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1176), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1169), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g764(.A(G319), .B1(new_n661), .B2(new_n662), .ZN(new_n1191));
  OR3_X1    g765(.A1(G227), .A2(KEYINPUT127), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g766(.A(KEYINPUT127), .B1(G227), .B2(new_n1191), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n703), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n1194), .A2(new_n921), .A3(new_n1003), .ZN(G225));
  INV_X1    g769(.A(G225), .ZN(G308));
endmodule


