//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT75), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  OR3_X1    g012(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n207), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n213), .ZN(new_n219));
  INV_X1    g018(.A(new_n205), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT29), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G197gat), .B(G204gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  INV_X1    g026(.A(G211gat), .ZN(new_n228));
  INV_X1    g027(.A(G218gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G211gat), .B(G218gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n226), .A3(new_n230), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT80), .B1(new_n225), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n207), .A2(new_n212), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n213), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n221), .ZN(new_n241));
  INV_X1    g040(.A(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n224), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247));
  INV_X1    g046(.A(new_n236), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G228gat), .A2(G233gat), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n234), .A2(KEYINPUT79), .A3(new_n235), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n231), .A2(new_n252), .A3(new_n233), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n245), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n224), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n237), .A2(new_n249), .A3(new_n250), .A4(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n225), .A2(new_n236), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n245), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n223), .B1(new_n260), .B2(new_n224), .ZN(new_n261));
  OAI211_X1 g060(.A(G228gat), .B(G233gat), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n258), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n258), .B2(new_n262), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n204), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n258), .A2(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n262), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n203), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273));
  INV_X1    g072(.A(G127gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n274), .B2(G134gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G113gat), .B(G120gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n277));
  XOR2_X1   g076(.A(G127gat), .B(G134gat), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G120gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G113gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n278), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n273), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n278), .A3(new_n275), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT76), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n291), .A3(new_n256), .ZN(new_n292));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n240), .A2(new_n243), .A3(new_n289), .A4(new_n290), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT39), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(new_n215), .B2(new_n222), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n244), .A2(new_n288), .A3(new_n299), .A4(new_n291), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n280), .A2(new_n287), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(new_n223), .A3(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n293), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT0), .ZN(new_n310));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n302), .A2(new_n304), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n293), .B1(new_n313), .B2(new_n300), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n314), .B2(new_n298), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT40), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n313), .A2(new_n319), .A3(new_n293), .A4(new_n300), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n300), .A2(new_n293), .A3(new_n302), .A4(new_n304), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT77), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT5), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n292), .A2(new_n294), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n306), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  OR3_X1    g125(.A1(new_n321), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT78), .B1(new_n321), .B2(KEYINPUT5), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n312), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n308), .A2(KEYINPUT40), .A3(new_n315), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n318), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G8gat), .B(G36gat), .Z(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G226gat), .ZN(new_n336));
  INV_X1    g135(.A(G233gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n341), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(KEYINPUT68), .A3(new_n347), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT27), .B(G183gat), .ZN(new_n352));
  INV_X1    g151(.A(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT28), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n350), .A2(new_n351), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(new_n340), .B2(KEYINPUT23), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n362), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n365));
  INV_X1    g164(.A(G176gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n365), .A2(KEYINPUT23), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n343), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n372), .A2(new_n373), .B1(new_n347), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n359), .B1(new_n369), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT25), .A3(new_n343), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n361), .B2(new_n363), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n374), .A2(new_n347), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n370), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n358), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n338), .B1(new_n384), .B2(new_n245), .ZN(new_n385));
  AOI211_X1 g184(.A(new_n336), .B(new_n337), .C1(new_n358), .C2(new_n383), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n248), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n338), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n358), .B2(new_n383), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n388), .B(new_n236), .C1(new_n338), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n335), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n390), .A3(new_n335), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n387), .A2(KEYINPUT30), .A3(new_n390), .A4(new_n335), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n272), .B1(new_n332), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n387), .A2(new_n390), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT37), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT37), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n387), .A2(KEYINPUT82), .A3(new_n390), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT38), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n335), .B1(new_n402), .B2(KEYINPUT37), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n329), .A2(KEYINPUT6), .A3(new_n312), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  INV_X1    g210(.A(new_n312), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n326), .A2(new_n327), .A3(new_n412), .A4(new_n328), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n330), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n409), .A2(new_n410), .A3(new_n414), .A4(new_n393), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n400), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n358), .A2(new_n383), .A3(new_n303), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n303), .B1(new_n358), .B2(new_n383), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G71gat), .B(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n433));
  INV_X1    g232(.A(new_n303), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n372), .A2(new_n373), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n380), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n368), .A2(new_n343), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n364), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n438), .A2(new_n359), .B1(new_n381), .B2(new_n379), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n346), .A2(KEYINPUT68), .A3(new_n347), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT68), .B1(new_n346), .B2(new_n347), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n355), .A2(new_n357), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n434), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n421), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n433), .B1(new_n445), .B2(new_n420), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n426), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT70), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AND4_X1   g248(.A1(KEYINPUT70), .A2(new_n424), .A3(KEYINPUT32), .A4(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n432), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n445), .A2(new_n420), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n452), .B(new_n453), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n432), .C1(new_n449), .C2(new_n450), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT72), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n451), .A2(new_n454), .A3(KEYINPUT72), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT36), .ZN(new_n463));
  INV_X1    g262(.A(new_n399), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n414), .A2(new_n410), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n462), .A2(new_n463), .B1(new_n466), .B2(new_n272), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n400), .B(KEYINPUT83), .C1(new_n415), .C2(new_n416), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n419), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n267), .A2(new_n271), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n457), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT84), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n399), .B1(new_n410), .B2(new_n414), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n470), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n461), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n272), .A2(KEYINPUT35), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n473), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n469), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT87), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G8gat), .ZN(new_n485));
  INV_X1    g284(.A(G8gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(KEYINPUT87), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  AOI21_X1  g288(.A(G1gat), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n490), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(G71gat), .A2(G78gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(G71gat), .A2(G78gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n499), .ZN(new_n502));
  INV_X1    g301(.A(G57gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G64gat), .ZN(new_n504));
  INV_X1    g303(.A(G64gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G57gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n501), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT21), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT90), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n513), .B(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n509), .A2(KEYINPUT21), .ZN(new_n519));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G183gat), .B(G211gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n518), .B(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G43gat), .ZN(new_n529));
  INV_X1    g328(.A(G50gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G43gat), .A2(G50gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT85), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(KEYINPUT15), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535));
  INV_X1    g334(.A(G29gat), .ZN(new_n536));
  INV_X1    g335(.A(G36gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT14), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G29gat), .B2(G36gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT86), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n535), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n542), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n534), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n528), .A2(KEYINPUT15), .A3(new_n533), .ZN(new_n547));
  INV_X1    g346(.A(new_n541), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n549), .A3(new_n532), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n535), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n525), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n545), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n547), .B1(new_n554), .B2(new_n543), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n548), .A3(new_n535), .A4(new_n550), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT17), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n559), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n563), .B2(new_n564), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n568), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n557), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT92), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n555), .A2(new_n556), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n583), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n579), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n582), .ZN(new_n592));
  XOR2_X1   g391(.A(G134gat), .B(G162gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n578), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n589), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n597), .A2(KEYINPUT93), .A3(new_n589), .A4(new_n594), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n524), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n507), .A2(new_n501), .A3(new_n502), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n607), .A3(KEYINPUT95), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n576), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n605), .B(new_n606), .C1(new_n585), .C2(new_n586), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n575), .B(new_n570), .C1(new_n500), .C2(new_n508), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n604), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n616), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n604), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(KEYINPUT96), .B(new_n604), .C1(new_n612), .C2(new_n617), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n625), .B1(new_n629), .B2(new_n624), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n603), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n553), .A2(new_n494), .A3(new_n557), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT88), .Z(new_n635));
  INV_X1    g434(.A(new_n494), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n584), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT18), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n635), .B(KEYINPUT13), .Z(new_n641));
  NOR2_X1   g440(.A1(new_n636), .A2(new_n584), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n494), .B1(new_n555), .B2(new_n556), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n633), .A2(KEYINPUT18), .A3(new_n637), .A4(new_n635), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT12), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n640), .A2(new_n644), .A3(new_n645), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT89), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n649), .B(KEYINPUT12), .Z(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n638), .B2(new_n639), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT89), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n644), .A4(new_n645), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n644), .A3(new_n645), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n632), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n482), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n465), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g465(.A(new_n486), .B1(new_n663), .B2(new_n399), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n662), .A2(new_n464), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  NAND2_X1  g470(.A1(new_n462), .A2(new_n463), .ZN(new_n672));
  OAI21_X1  g471(.A(G15gat), .B1(new_n662), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(G15gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n478), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n662), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT98), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n470), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n482), .A2(new_n601), .ZN(new_n681));
  INV_X1    g480(.A(new_n660), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(new_n524), .A3(new_n630), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n536), .A3(new_n664), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n482), .A2(KEYINPUT99), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n469), .A2(new_n481), .A3(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n602), .A2(KEYINPUT44), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n683), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n465), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n687), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n685), .A2(new_n537), .A3(new_n399), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n464), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n478), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n529), .ZN(new_n703));
  INV_X1    g502(.A(new_n672), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G43gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT100), .B(KEYINPUT47), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n706), .B(new_n707), .Z(G1330gat));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n681), .A2(G50gat), .A3(new_n470), .A4(new_n684), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n272), .A3(new_n683), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(G50gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n684), .B1(new_n692), .B2(new_n693), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n530), .B1(new_n715), .B2(new_n272), .ZN(new_n716));
  OAI211_X1 g515(.A(KEYINPUT101), .B(KEYINPUT48), .C1(new_n716), .C2(new_n710), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n714), .A2(new_n717), .ZN(G1331gat));
  INV_X1    g517(.A(new_n630), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n603), .A2(new_n660), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n688), .A2(new_n690), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT102), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n688), .A2(new_n723), .A3(new_n690), .A4(new_n720), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n664), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g525(.A(new_n464), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n729), .B(new_n730), .Z(G1333gat));
  XNOR2_X1  g530(.A(new_n478), .B(KEYINPUT104), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n722), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(G71gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n722), .A2(G71gat), .A3(new_n704), .A4(new_n724), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n272), .A3(new_n724), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT105), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n660), .A2(new_n524), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n719), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n694), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n465), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n681), .B2(new_n743), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n482), .A2(KEYINPUT51), .A3(new_n601), .A4(new_n742), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT106), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n664), .A2(new_n563), .A3(new_n630), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n746), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n694), .A2(new_n399), .A3(new_n744), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(new_n749), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n464), .A2(G92gat), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(new_n630), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n564), .B1(new_n755), .B2(KEYINPUT107), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n694), .A2(new_n762), .A3(new_n399), .A4(new_n744), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n759), .A2(KEYINPUT52), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(G1337gat));
  XNOR2_X1  g565(.A(KEYINPUT108), .B(G99gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n478), .A2(new_n630), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n745), .A2(new_n672), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n752), .A2(new_n768), .B1(new_n769), .B2(new_n767), .ZN(G1338gat));
  INV_X1    g569(.A(new_n744), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n470), .B(new_n771), .C1(new_n692), .C2(new_n693), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT109), .B(G106gat), .Z(new_n773));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n470), .A2(G106gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n630), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n772), .B2(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI221_X1 g578(.A(new_n776), .B1(KEYINPUT110), .B2(KEYINPUT53), .C1(new_n772), .C2(new_n773), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1339gat));
  INV_X1    g580(.A(new_n524), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n612), .A2(new_n617), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(new_n604), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n618), .A2(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n627), .A2(new_n789), .A3(new_n628), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791));
  INV_X1    g590(.A(new_n624), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n791), .B1(new_n790), .B2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n788), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n787), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n790), .A2(new_n792), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT111), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(new_n793), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n625), .B(new_n796), .C1(new_n801), .C2(KEYINPUT55), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n642), .A2(new_n643), .A3(new_n641), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n635), .B1(new_n633), .B2(new_n637), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n649), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n657), .A2(new_n601), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n783), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n657), .A2(new_n601), .A3(new_n805), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n797), .B1(new_n794), .B2(new_n795), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n784), .ZN(new_n810));
  INV_X1    g609(.A(new_n625), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n800), .A2(new_n793), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n788), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(KEYINPUT112), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n810), .A2(new_n813), .A3(new_n660), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n657), .A2(new_n630), .A3(new_n805), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n601), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n782), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n682), .A2(new_n602), .A3(new_n524), .A4(new_n719), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT113), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n472), .A2(new_n475), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n399), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n825), .A2(new_n664), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n282), .A3(new_n660), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n465), .A2(new_n399), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n478), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n823), .B1(new_n819), .B2(new_n820), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n470), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n470), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n833), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n660), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n831), .B1(new_n841), .B2(G113gat), .ZN(new_n842));
  AOI211_X1 g641(.A(KEYINPUT115), .B(new_n282), .C1(new_n840), .C2(new_n660), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n830), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  AOI21_X1  g643(.A(G120gat), .B1(new_n829), .B2(new_n630), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n719), .A2(new_n284), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n840), .B2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(new_n833), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n782), .A2(new_n274), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n838), .B1(new_n825), .B2(new_n470), .ZN(new_n850));
  INV_X1    g649(.A(new_n839), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n840), .A2(KEYINPUT116), .A3(new_n849), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n274), .B1(new_n828), .B2(new_n782), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT117), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n854), .A2(new_n855), .A3(new_n859), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1342gat));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n602), .A2(G134gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n829), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n863), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT56), .B1(new_n828), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n840), .A2(new_n601), .ZN(new_n868));
  INV_X1    g667(.A(G134gat), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n867), .B(KEYINPUT118), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n840), .B2(new_n601), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n864), .A2(new_n866), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(G1343gat));
  NAND2_X1  g674(.A1(new_n672), .A2(new_n832), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n825), .B2(new_n272), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n272), .A2(KEYINPUT57), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n819), .B2(new_n820), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n660), .B(new_n877), .C1(new_n878), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT58), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n660), .A2(new_n208), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n704), .A2(new_n470), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n664), .B(new_n885), .C1(new_n834), .C2(new_n835), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT119), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n825), .A2(new_n888), .A3(new_n664), .A4(new_n885), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n889), .A3(new_n464), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n886), .A2(new_n399), .A3(new_n884), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n882), .B2(G141gat), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1344gat));
  OAI21_X1  g694(.A(KEYINPUT59), .B1(new_n890), .B2(new_n719), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n209), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n877), .B1(new_n878), .B2(new_n881), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n719), .A2(KEYINPUT59), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n632), .A2(new_n682), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n802), .A2(new_n806), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n782), .B1(new_n818), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n470), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(KEYINPUT120), .A3(new_n903), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n880), .B1(new_n822), .B2(new_n824), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n719), .A3(new_n876), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n897), .B(new_n900), .C1(new_n911), .C2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n898), .B2(new_n782), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n524), .A2(new_n216), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n890), .B2(new_n915), .ZN(G1346gat));
  OAI21_X1  g715(.A(new_n217), .B1(new_n890), .B2(new_n602), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n602), .A2(new_n217), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n877), .B(new_n918), .C1(new_n878), .C2(new_n881), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n826), .A2(new_n464), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n465), .B1(new_n834), .B2(new_n835), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n825), .A2(new_n929), .A3(new_n465), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n931), .A2(new_n365), .A3(new_n367), .A4(new_n660), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n664), .A2(new_n464), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n732), .A2(new_n933), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n682), .B(new_n934), .C1(new_n837), .C2(new_n839), .ZN(new_n935));
  INV_X1    g734(.A(G169gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  NAND2_X1  g736(.A1(new_n837), .A2(new_n839), .ZN(new_n938));
  INV_X1    g737(.A(new_n934), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n719), .A2(new_n366), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n938), .A2(KEYINPUT124), .A3(new_n939), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n931), .A2(new_n630), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT123), .B1(new_n946), .B2(new_n366), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n948), .B(G176gat), .C1(new_n931), .C2(new_n630), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(G1349gat));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n524), .A2(new_n352), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n931), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n524), .B(new_n939), .C1(new_n850), .C2(new_n851), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G183gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n951), .A2(new_n952), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n955), .B2(new_n957), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n931), .A2(new_n353), .A3(new_n601), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n938), .A2(new_n601), .A3(new_n939), .ZN(new_n963));
  XNOR2_X1  g762(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(G190gat), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n963), .B2(G190gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1351gat));
  NAND2_X1  g766(.A1(new_n672), .A2(new_n933), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n910), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n682), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n928), .A2(new_n930), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n704), .A2(new_n464), .A3(new_n470), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n660), .A3(new_n973), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n969), .A2(new_n971), .B1(new_n970), .B2(new_n974), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n719), .A2(G204gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n977), .A2(KEYINPUT62), .ZN(new_n979));
  INV_X1    g778(.A(new_n968), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n630), .B(new_n980), .C1(new_n908), .C2(new_n909), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n981), .A2(KEYINPUT127), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n978), .B(new_n979), .C1(new_n983), .C2(new_n984), .ZN(G1353gat));
  OAI211_X1 g784(.A(new_n524), .B(new_n980), .C1(new_n908), .C2(new_n909), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n524), .A2(new_n228), .ZN(new_n990));
  OAI22_X1  g789(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n990), .ZN(G1354gat));
  AOI21_X1  g790(.A(new_n229), .B1(new_n969), .B2(new_n601), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n989), .A2(G218gat), .A3(new_n602), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n992), .A2(new_n993), .ZN(G1355gat));
endmodule


