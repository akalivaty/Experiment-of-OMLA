

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n457), .B(n456), .Z(n290) );
  XNOR2_X1 U323 ( .A(n291), .B(n392), .ZN(n394) );
  XOR2_X1 U324 ( .A(n476), .B(KEYINPUT28), .Z(n525) );
  XOR2_X1 U325 ( .A(n437), .B(n387), .Z(n291) );
  INV_X1 U326 ( .A(KEYINPUT25), .ZN(n404) );
  XNOR2_X1 U327 ( .A(n404), .B(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U328 ( .A(n406), .B(n405), .ZN(n410) );
  INV_X1 U329 ( .A(KEYINPUT115), .ZN(n459) );
  XNOR2_X1 U330 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U331 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n470) );
  INV_X1 U332 ( .A(KEYINPUT23), .ZN(n396) );
  XNOR2_X1 U333 ( .A(n471), .B(n470), .ZN(n531) );
  XNOR2_X1 U334 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U335 ( .A(n416), .B(KEYINPUT100), .ZN(n417) );
  XNOR2_X1 U336 ( .A(n399), .B(n398), .ZN(n400) );
  NOR2_X1 U337 ( .A1(n475), .A2(n517), .ZN(n570) );
  XNOR2_X1 U338 ( .A(n418), .B(n417), .ZN(n516) );
  XOR2_X1 U339 ( .A(KEYINPUT18), .B(n346), .Z(n384) );
  XOR2_X1 U340 ( .A(n461), .B(KEYINPUT81), .Z(n543) );
  XOR2_X1 U341 ( .A(n384), .B(n383), .Z(n522) );
  XNOR2_X1 U342 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U343 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U344 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n454), .B(n453), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G71GAT), .Z(n293) );
  XNOR2_X1 U347 ( .A(G183GAT), .B(G127GAT), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U349 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n295) );
  XNOR2_X1 U350 ( .A(G8GAT), .B(KEYINPUT82), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n434) );
  XOR2_X1 U354 ( .A(G155GAT), .B(G78GAT), .Z(n299) );
  XNOR2_X1 U355 ( .A(G22GAT), .B(G211GAT), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n434), .B(n300), .Z(n302) );
  NAND2_X1 U358 ( .A1(G231GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U360 ( .A(n303), .B(KEYINPUT15), .Z(n306) );
  XNOR2_X1 U361 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n304), .B(KEYINPUT71), .ZN(n426) );
  XNOR2_X1 U363 ( .A(n426), .B(KEYINPUT83), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U365 ( .A(n308), .B(n307), .Z(n567) );
  INV_X1 U366 ( .A(n567), .ZN(n578) );
  INV_X1 U367 ( .A(KEYINPUT36), .ZN(n331) );
  XOR2_X1 U368 ( .A(G43GAT), .B(G29GAT), .Z(n310) );
  XNOR2_X1 U369 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U371 ( .A(n311), .B(KEYINPUT68), .Z(n313) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n448) );
  XOR2_X1 U374 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U377 ( .A(KEYINPUT10), .B(KEYINPUT64), .Z(n317) );
  XNOR2_X1 U378 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n329) );
  XOR2_X1 U381 ( .A(KEYINPUT76), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U382 ( .A(G190GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n320), .B(KEYINPUT79), .ZN(n341) );
  XNOR2_X1 U384 ( .A(n387), .B(n341), .ZN(n322) );
  AND2_X1 U385 ( .A1(G232GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U387 ( .A(KEYINPUT74), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U390 ( .A(G106GAT), .B(KEYINPUT73), .Z(n325) );
  XOR2_X1 U391 ( .A(n326), .B(n325), .Z(n430) );
  XNOR2_X1 U392 ( .A(n327), .B(n430), .ZN(n328) );
  XOR2_X1 U393 ( .A(n329), .B(n328), .Z(n330) );
  XNOR2_X1 U394 ( .A(n448), .B(n330), .ZN(n461) );
  XNOR2_X1 U395 ( .A(n331), .B(n543), .ZN(n455) );
  XOR2_X1 U396 ( .A(G64GAT), .B(KEYINPUT75), .Z(n333) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n427) );
  XOR2_X1 U399 ( .A(G169GAT), .B(G8GAT), .Z(n433) );
  XOR2_X1 U400 ( .A(n427), .B(n433), .Z(n335) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U403 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n337) );
  XNOR2_X1 U404 ( .A(G36GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U405 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U406 ( .A(n339), .B(n338), .Z(n343) );
  XNOR2_X1 U407 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n340), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U409 ( .A(n386), .B(n341), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U411 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n345) );
  XNOR2_X1 U412 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U414 ( .A(n347), .B(n384), .Z(n472) );
  INV_X1 U415 ( .A(n472), .ZN(n520) );
  XNOR2_X1 U416 ( .A(n520), .B(KEYINPUT27), .ZN(n408) );
  XOR2_X1 U417 ( .A(G148GAT), .B(G120GAT), .Z(n349) );
  XNOR2_X1 U418 ( .A(G29GAT), .B(G141GAT), .ZN(n348) );
  XNOR2_X1 U419 ( .A(n349), .B(n348), .ZN(n351) );
  XOR2_X1 U420 ( .A(G162GAT), .B(G85GAT), .Z(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n360) );
  XOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n358) );
  XNOR2_X1 U423 ( .A(G127GAT), .B(KEYINPUT84), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n352), .B(KEYINPUT0), .ZN(n353) );
  XOR2_X1 U425 ( .A(n353), .B(KEYINPUT85), .Z(n355) );
  XNOR2_X1 U426 ( .A(G113GAT), .B(G134GAT), .ZN(n354) );
  XNOR2_X1 U427 ( .A(n355), .B(n354), .ZN(n380) );
  XNOR2_X1 U428 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n356) );
  XNOR2_X1 U429 ( .A(n356), .B(KEYINPUT2), .ZN(n395) );
  XNOR2_X1 U430 ( .A(n380), .B(n395), .ZN(n357) );
  XNOR2_X1 U431 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n360), .B(n359), .ZN(n362) );
  NAND2_X1 U433 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n370) );
  XOR2_X1 U435 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n364) );
  XNOR2_X1 U436 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n363) );
  XNOR2_X1 U437 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U438 ( .A(KEYINPUT90), .B(KEYINPUT93), .Z(n366) );
  XNOR2_X1 U439 ( .A(G1GAT), .B(G57GAT), .ZN(n365) );
  XNOR2_X1 U440 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U441 ( .A(n368), .B(n367), .Z(n369) );
  XNOR2_X1 U442 ( .A(n370), .B(n369), .ZN(n517) );
  NAND2_X1 U443 ( .A1(n408), .A2(n517), .ZN(n530) );
  XOR2_X1 U444 ( .A(G190GAT), .B(G99GAT), .Z(n372) );
  XNOR2_X1 U445 ( .A(G43GAT), .B(G15GAT), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U447 ( .A(n373), .B(KEYINPUT87), .Z(n375) );
  XOR2_X1 U448 ( .A(G120GAT), .B(G71GAT), .Z(n422) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(n422), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n377) );
  NAND2_X1 U452 ( .A1(G227GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U453 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U454 ( .A(n379), .B(n378), .Z(n382) );
  XNOR2_X1 U455 ( .A(n380), .B(G176GAT), .ZN(n381) );
  XNOR2_X1 U456 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U457 ( .A(n522), .ZN(n535) );
  XNOR2_X1 U458 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n385) );
  XNOR2_X1 U459 ( .A(n385), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U460 ( .A(n386), .B(n419), .ZN(n401) );
  XOR2_X1 U461 ( .A(G141GAT), .B(G22GAT), .Z(n437) );
  XOR2_X1 U462 ( .A(G106GAT), .B(G218GAT), .Z(n391) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n389) );
  XNOR2_X1 U464 ( .A(G50GAT), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U465 ( .A(n389), .B(n388), .ZN(n390) );
  NAND2_X1 U466 ( .A1(G228GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U467 ( .A(n394), .B(n393), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n395), .B(KEYINPUT22), .ZN(n397) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n476) );
  INV_X1 U470 ( .A(n525), .ZN(n533) );
  NAND2_X1 U471 ( .A1(n535), .A2(n533), .ZN(n402) );
  NOR2_X1 U472 ( .A1(n530), .A2(n402), .ZN(n414) );
  NAND2_X1 U473 ( .A1(n520), .A2(n522), .ZN(n403) );
  NAND2_X1 U474 ( .A1(n403), .A2(n476), .ZN(n406) );
  NOR2_X1 U475 ( .A1(n476), .A2(n522), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT26), .ZN(n569) );
  NAND2_X1 U477 ( .A1(n408), .A2(n569), .ZN(n409) );
  NAND2_X1 U478 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U479 ( .A(KEYINPUT97), .B(n411), .ZN(n412) );
  NOR2_X1 U480 ( .A1(n517), .A2(n412), .ZN(n413) );
  NOR2_X1 U481 ( .A1(n414), .A2(n413), .ZN(n485) );
  NOR2_X1 U482 ( .A1(n455), .A2(n485), .ZN(n415) );
  NAND2_X1 U483 ( .A1(n578), .A2(n415), .ZN(n418) );
  XNOR2_X1 U484 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n416) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(n419), .Z(n421) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n422), .B(KEYINPUT33), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n423), .B(KEYINPUT31), .ZN(n424) );
  XOR2_X1 U490 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U491 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n432) );
  XOR2_X1 U494 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U497 ( .A(n438), .B(n437), .Z(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n440) );
  XNOR2_X1 U499 ( .A(G197GAT), .B(G113GAT), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U501 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n442) );
  XNOR2_X1 U502 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n571) );
  XOR2_X1 U507 ( .A(n571), .B(KEYINPUT70), .Z(n559) );
  NAND2_X1 U508 ( .A1(n432), .A2(n559), .ZN(n488) );
  NOR2_X1 U509 ( .A1(n516), .A2(n488), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n449), .B(KEYINPUT102), .ZN(n450) );
  XNOR2_X1 U511 ( .A(KEYINPUT38), .B(n450), .ZN(n502) );
  NAND2_X1 U512 ( .A1(n502), .A2(n522), .ZN(n454) );
  XOR2_X1 U513 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n452) );
  XNOR2_X1 U514 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n451) );
  INV_X1 U515 ( .A(KEYINPUT54), .ZN(n474) );
  XOR2_X1 U516 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n457) );
  NOR2_X1 U517 ( .A1(n455), .A2(n578), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n432), .A2(n290), .ZN(n458) );
  NOR2_X1 U519 ( .A1(n458), .A2(n559), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n469) );
  INV_X1 U521 ( .A(KEYINPUT47), .ZN(n467) );
  XOR2_X1 U522 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n463) );
  XOR2_X1 U523 ( .A(KEYINPUT41), .B(n432), .Z(n550) );
  NOR2_X1 U524 ( .A1(n571), .A2(n550), .ZN(n462) );
  XOR2_X1 U525 ( .A(n463), .B(n462), .Z(n464) );
  NAND2_X1 U526 ( .A1(n578), .A2(n464), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n461), .A2(n465), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n531), .A2(n472), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n570), .A2(n476), .ZN(n478) );
  XOR2_X1 U533 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X2 U535 ( .A1(n479), .A2(n535), .ZN(n566) );
  NAND2_X1 U536 ( .A1(n566), .A2(n543), .ZN(n483) );
  XOR2_X1 U537 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n481) );
  INV_X1 U538 ( .A(G190GAT), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n578), .A2(n543), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n484), .B(KEYINPUT16), .ZN(n487) );
  INV_X1 U541 ( .A(n485), .ZN(n486) );
  NAND2_X1 U542 ( .A1(n487), .A2(n486), .ZN(n505) );
  NOR2_X1 U543 ( .A1(n488), .A2(n505), .ZN(n496) );
  NAND2_X1 U544 ( .A1(n517), .A2(n496), .ZN(n491) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT98), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n520), .A2(n496), .ZN(n492) );
  XNOR2_X1 U549 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U551 ( .A1(n496), .A2(n522), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n495), .Z(G1326GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n525), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U557 ( .A1(n502), .A2(n517), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT103), .Z(n501) );
  NAND2_X1 U560 ( .A1(n502), .A2(n520), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n504) );
  NAND2_X1 U563 ( .A1(n525), .A2(n502), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n550), .B(KEYINPUT107), .ZN(n561) );
  NAND2_X1 U567 ( .A1(n571), .A2(n561), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n515), .A2(n505), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n512), .A2(n517), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n520), .A2(n512), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(KEYINPUT108), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U575 ( .A1(n512), .A2(n522), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U578 ( .A1(n512), .A2(n525), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n519) );
  NOR2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n526), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT111), .Z(n524) );
  NAND2_X1 U587 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n528) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT117), .B(n532), .Z(n548) );
  NAND2_X1 U595 ( .A1(n548), .A2(n533), .ZN(n534) );
  NOR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n559), .A2(n544), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(KEYINPUT118), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n544), .A2(n561), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n541) );
  NAND2_X1 U604 ( .A1(n544), .A2(n567), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n548), .A2(n569), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n571), .A2(n556), .ZN(n549) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n556), .A2(n550), .ZN(n554) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n578), .A2(n556), .ZN(n555) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  INV_X1 U621 ( .A(n556), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n557), .A2(n461), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n566), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n566), .A2(n561), .ZN(n563) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n581), .A2(n571), .ZN(n575) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n573) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n432), .A2(n581), .ZN(n577) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n581), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n455), .A2(n581), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

