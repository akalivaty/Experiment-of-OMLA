//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n209), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT14), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT15), .A3(new_n213), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n214), .A2(new_n218), .A3(new_n222), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT88), .A2(KEYINPUT17), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT88), .A2(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n212), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n212), .A2(new_n224), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n234), .A2(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(KEYINPUT18), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n231), .B(KEYINPUT13), .Z(new_n237));
  NOR2_X1   g036(.A1(new_n212), .A2(new_n224), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT11), .ZN(new_n242));
  INV_X1    g041(.A(G169gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT89), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n235), .A2(new_n246), .A3(new_n236), .A4(new_n239), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n248), .B2(new_n250), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G57gat), .B(G85gat), .Z(new_n255));
  XNOR2_X1  g054(.A(G1gat), .B(G29gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n257), .B(new_n258), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n260));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT76), .A2(G148gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(G141gat), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G148gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n264), .A2(new_n266), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n270), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n267), .ZN(new_n274));
  XOR2_X1   g073(.A(G141gat), .B(G148gat), .Z(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(new_n268), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G127gat), .B(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g079(.A1(G113gat), .A2(G120gat), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n279), .A2(new_n280), .A3(new_n281), .A4(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n280), .A3(new_n281), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(G113gat), .B2(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n281), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT68), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(new_n290), .A3(new_n278), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n277), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(new_n277), .B2(new_n292), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n261), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n275), .A2(new_n268), .ZN(new_n299));
  INV_X1    g098(.A(new_n274), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n264), .A2(new_n266), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n271), .A2(new_n267), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n291), .A3(KEYINPUT77), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(new_n272), .B2(new_n276), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n298), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n260), .B1(new_n296), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g110(.A(new_n277), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(new_n312), .A3(new_n306), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n277), .A2(new_n292), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n261), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(KEYINPUT4), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n277), .A2(new_n292), .A3(new_n293), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT78), .A3(new_n308), .A4(new_n261), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n310), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n318), .A2(KEYINPUT80), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(new_n309), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n318), .A2(KEYINPUT80), .A3(new_n319), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(new_n311), .A3(new_n261), .A4(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n259), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT6), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(KEYINPUT81), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT6), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n326), .A3(new_n259), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n331), .B(new_n332), .C1(new_n327), .C2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337));
  INV_X1    g136(.A(G211gat), .ZN(new_n338));
  INV_X1    g137(.A(G218gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n336), .A3(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  INV_X1    g148(.A(G176gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n243), .A2(new_n350), .A3(KEYINPUT23), .ZN(new_n351));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n351), .A2(KEYINPUT65), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT65), .B1(new_n351), .B2(new_n352), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G190gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(G183gat), .ZN(new_n357));
  INV_X1    g156(.A(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G190gat), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(KEYINPUT24), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n243), .A2(new_n350), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n360), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n349), .B1(new_n355), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n352), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n365), .B2(new_n366), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(KEYINPUT23), .A3(new_n243), .A4(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n360), .A2(new_n371), .A3(new_n363), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n364), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT65), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n366), .A2(G169gat), .A3(G176gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(new_n370), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n351), .A2(KEYINPUT65), .A3(new_n352), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n358), .A2(G190gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n356), .A2(G183gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n362), .B1(new_n384), .B2(KEYINPUT24), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n381), .A2(KEYINPUT66), .A3(new_n385), .A4(new_n367), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n376), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT27), .B(G183gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n356), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT28), .B1(new_n389), .B2(KEYINPUT67), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n391), .B(new_n392), .C1(new_n388), .C2(new_n356), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n352), .B1(new_n365), .B2(KEYINPUT26), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n361), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OR3_X1    g196(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(G226gat), .ZN(new_n400));
  INV_X1    g199(.A(G233gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n348), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n385), .B(new_n367), .C1(new_n354), .C2(new_n353), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(new_n349), .B1(new_n364), .B2(new_n375), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n386), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT72), .B(new_n404), .C1(new_n408), .C2(KEYINPUT29), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n387), .A2(new_n398), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT73), .B1(new_n411), .B2(new_n402), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n413), .B(new_n404), .C1(new_n387), .C2(new_n398), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n347), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G64gat), .ZN(new_n418));
  INV_X1    g217(.A(G92gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n402), .B1(new_n411), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n404), .B1(new_n387), .B2(new_n398), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n422), .A2(new_n347), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT30), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n416), .A2(new_n425), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT74), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n416), .A2(new_n430), .A3(new_n425), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n420), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT75), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n403), .B(new_n409), .C1(new_n412), .C2(new_n414), .ZN(new_n435));
  AOI211_X1 g234(.A(KEYINPUT74), .B(new_n424), .C1(new_n435), .C2(new_n347), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n416), .B2(new_n425), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT75), .B(new_n433), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n335), .B(new_n427), .C1(new_n434), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n346), .A2(new_n421), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n302), .B1(new_n442), .B2(KEYINPUT83), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT29), .B1(new_n344), .B2(new_n345), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT83), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n312), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n277), .B2(new_n302), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n346), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n441), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n312), .B(new_n452), .C1(KEYINPUT3), .C2(new_n444), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT82), .B(new_n307), .C1(new_n442), .C2(new_n277), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n441), .B1(new_n448), .B2(new_n346), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(G22gat), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n450), .A2(new_n454), .A3(new_n441), .A4(new_n453), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT3), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n277), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(G228gat), .B(G233gat), .C1(new_n462), .C2(new_n449), .ZN(new_n463));
  INV_X1    g262(.A(G22gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT31), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n467), .B(G50gat), .Z(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT84), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n458), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n458), .B2(new_n465), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n411), .A2(new_n292), .ZN(new_n475));
  INV_X1    g274(.A(G227gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n401), .ZN(new_n477));
  INV_X1    g276(.A(new_n292), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n387), .A2(new_n478), .A3(new_n398), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(G71gat), .B(G99gat), .Z(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n480), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n480), .A2(new_n484), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n483), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n477), .B1(new_n475), .B2(new_n479), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  INV_X1    g298(.A(new_n479), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n478), .B1(new_n387), .B2(new_n398), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n500), .A2(new_n501), .B1(new_n476), .B2(new_n401), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n502), .B2(KEYINPUT71), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n491), .A3(new_n494), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n474), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT35), .B1(new_n440), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n427), .B1(new_n434), .B2(new_n439), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n513));
  AND3_X1   g312(.A1(new_n504), .A2(new_n491), .A3(new_n494), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n504), .B1(new_n491), .B2(new_n494), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n470), .B2(new_n473), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n328), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n506), .A2(KEYINPUT85), .A3(new_n507), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n511), .B1(new_n512), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n516), .A2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n426), .B(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n529), .B2(new_n438), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(new_n530), .A3(KEYINPUT86), .A4(new_n520), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n523), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n332), .A2(new_n331), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n328), .B(new_n426), .C1(new_n533), .C2(new_n327), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n428), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n422), .ZN(new_n537));
  INV_X1    g336(.A(new_n423), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n347), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n347), .B2(new_n435), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n420), .A2(KEYINPUT38), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n534), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n429), .A2(KEYINPUT37), .A3(new_n431), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n420), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n474), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n261), .B1(new_n324), .B2(new_n325), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT39), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT39), .B1(new_n315), .B2(new_n316), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n552), .B(new_n259), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n327), .B1(new_n555), .B2(KEYINPUT40), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(KEYINPUT40), .B2(new_n555), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n548), .B(new_n549), .C1(new_n530), .C2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n514), .B2(new_n515), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n506), .A2(KEYINPUT36), .A3(new_n507), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n440), .B2(new_n474), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n254), .B1(new_n532), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n572), .B2(new_n419), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  AOI21_X1  g375(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT90), .B1(new_n581), .B2(G57gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT90), .A3(G57gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(G57gat), .B2(new_n581), .ZN(new_n584));
  OAI221_X1 g383(.A(new_n580), .B1(new_n579), .B2(new_n578), .C1(new_n582), .C2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n588), .A2(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n568), .B1(new_n576), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n574), .B(new_n575), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(new_n589), .A3(new_n585), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT10), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n567), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n594), .A2(new_n567), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G176gat), .ZN(new_n602));
  INV_X1    g401(.A(G204gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n597), .B1(new_n594), .B2(new_n595), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT94), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n567), .B1(new_n607), .B2(KEYINPUT94), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n599), .B(new_n604), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n566), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n611), .A3(new_n566), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n228), .A2(new_n229), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n576), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n224), .A2(new_n592), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n618), .A2(new_n630), .A3(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n626), .B2(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n210), .B(new_n211), .C1(new_n590), .C2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n358), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT92), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n639), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n590), .A2(new_n637), .ZN(new_n645));
  XOR2_X1   g444(.A(G127gat), .B(G155gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n338), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n648), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n616), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n565), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n335), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n512), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT16), .B(G8gat), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT42), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(G8gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT96), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1325gat));
  INV_X1    g465(.A(new_n524), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n655), .A2(G15gat), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n656), .A2(new_n562), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(G15gat), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT97), .Z(G1326gat));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n549), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(new_n651), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n615), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n636), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT98), .Z(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(new_n565), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n215), .A3(new_n657), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n633), .B2(new_n634), .ZN(new_n683));
  INV_X1    g482(.A(new_n634), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n632), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g485(.A(KEYINPUT44), .B(new_n686), .C1(new_n532), .C2(new_n564), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n532), .A2(new_n564), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n636), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n691), .B2(KEYINPUT44), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n635), .B1(new_n532), .B2(new_n564), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(KEYINPUT99), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n688), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n248), .A2(new_n250), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n676), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT101), .B1(new_n700), .B2(new_n335), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G29gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n700), .A2(KEYINPUT101), .A3(new_n335), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n681), .B1(new_n702), .B2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n679), .A2(new_n216), .A3(new_n512), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  OAI21_X1  g505(.A(G36gat), .B1(new_n700), .B2(new_n530), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n679), .A2(new_n709), .A3(new_n524), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n691), .A2(new_n689), .A3(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT99), .B1(new_n693), .B2(new_n694), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n687), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n562), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n698), .ZN(new_n715));
  OAI211_X1 g514(.A(KEYINPUT47), .B(new_n710), .C1(new_n715), .C2(new_n709), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n715), .B2(new_n709), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT102), .B(G43gat), .C1(new_n700), .C2(new_n714), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n719), .A3(new_n710), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT103), .B1(new_n720), .B2(new_n721), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(G1330gat));
  NAND3_X1  g523(.A1(new_n696), .A2(new_n474), .A3(new_n699), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n549), .A2(G50gat), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n725), .A2(G50gat), .B1(new_n679), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g527(.A(new_n697), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n615), .A2(new_n729), .A3(new_n652), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n690), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n335), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT104), .B(G57gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n530), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(G1333gat));
  NOR3_X1   g538(.A1(new_n731), .A2(G71gat), .A3(new_n667), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n690), .A2(new_n562), .A3(new_n730), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(G71gat), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT105), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n731), .A2(new_n549), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(G78gat), .Z(G1335gat));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n691), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  AOI211_X1 g550(.A(new_n697), .B(new_n675), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n751), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n754), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n748), .A2(new_n756), .A3(new_n749), .A4(new_n752), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n615), .A2(new_n572), .A3(new_n657), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT109), .Z(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n696), .A2(new_n729), .A3(new_n651), .A4(new_n615), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n335), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1336gat));
  NOR2_X1   g565(.A1(new_n530), .A2(G92gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n758), .A2(new_n615), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n764), .A2(new_n530), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n419), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n769), .B2(new_n419), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI221_X1 g572(.A(new_n768), .B1(KEYINPUT110), .B2(KEYINPUT52), .C1(new_n769), .C2(new_n419), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1337gat));
  NOR3_X1   g574(.A1(new_n616), .A2(new_n667), .A3(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G99gat), .B1(new_n764), .B2(new_n714), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1338gat));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n549), .A2(G106gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n758), .A2(new_n615), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G106gat), .B1(new_n764), .B2(new_n549), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n784), .B(new_n786), .ZN(G1339gat));
  INV_X1    g586(.A(new_n686), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n607), .A2(KEYINPUT94), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n567), .A3(new_n608), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  INV_X1    g590(.A(new_n567), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n607), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n605), .B1(new_n598), .B2(KEYINPUT54), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT55), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(new_n697), .A3(new_n611), .A4(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n233), .A2(new_n238), .A3(new_n237), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT112), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n230), .A2(new_n233), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n231), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n245), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n250), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n614), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n612), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n788), .B1(new_n801), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n795), .B1(new_n790), .B2(new_n793), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n611), .B1(new_n812), .B2(KEYINPUT55), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT55), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n813), .A2(new_n814), .A3(new_n686), .A4(new_n807), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n651), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n654), .A2(new_n729), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n474), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n524), .B1(new_n818), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n512), .A2(new_n335), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n254), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n335), .B1(new_n816), .B2(new_n817), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n508), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n530), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n697), .A2(new_n282), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(KEYINPUT114), .Z(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n825), .A2(new_n831), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n824), .B2(new_n616), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n615), .A2(new_n283), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT115), .Z(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n824), .B2(new_n651), .ZN(new_n838));
  INV_X1    g637(.A(G127gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n828), .A2(new_n839), .A3(new_n675), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n512), .A2(new_n635), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT116), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n822), .A2(new_n636), .A3(new_n823), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n848), .A3(G134gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(G134gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n816), .A2(new_n817), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT119), .B(new_n854), .C1(new_n855), .C2(new_n549), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n653), .A2(new_n697), .ZN(new_n858));
  INV_X1    g657(.A(new_n815), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n813), .A2(new_n814), .ZN(new_n860));
  INV_X1    g659(.A(new_n253), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n251), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n860), .A2(new_n862), .B1(new_n615), .B2(new_n808), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n636), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n858), .B1(new_n864), .B2(new_n651), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n549), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n857), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n549), .B1(new_n816), .B2(new_n817), .ZN(new_n871));
  INV_X1    g670(.A(new_n854), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n799), .A2(new_n611), .A3(new_n800), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n810), .B1(new_n254), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n635), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n675), .B1(new_n876), .B2(new_n859), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT120), .B(new_n867), .C1(new_n877), .C2(new_n858), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n856), .A2(new_n869), .A3(new_n873), .A4(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n512), .A2(new_n562), .A3(new_n335), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n697), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G141gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n826), .A2(new_n474), .A3(new_n714), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n512), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n254), .A2(G141gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n853), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n853), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n879), .A2(new_n862), .A3(new_n880), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(G141gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n852), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(new_n888), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n881), .A2(G141gat), .B1(new_n884), .B2(new_n885), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n894), .B(KEYINPUT121), .C1(new_n853), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n891), .A2(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n880), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n616), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n262), .A2(new_n263), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n901), .A3(new_n615), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n880), .B(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n860), .A2(new_n636), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n807), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n876), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n912), .A2(new_n651), .B1(new_n254), .B2(new_n654), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n866), .B1(new_n913), .B2(new_n549), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n871), .A2(new_n872), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n616), .B(new_n907), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n917));
  OAI221_X1 g716(.A(new_n902), .B1(new_n905), .B2(new_n906), .C1(new_n916), .C2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n899), .B2(new_n651), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n884), .A2(new_n269), .A3(new_n675), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n899), .B2(new_n686), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n843), .A2(new_n270), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n883), .B2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n855), .A2(new_n657), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n512), .A3(new_n508), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n243), .A3(new_n697), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT125), .ZN(new_n929));
  INV_X1    g728(.A(new_n822), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n530), .A2(new_n657), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n930), .A2(new_n254), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n933), .B2(new_n243), .ZN(G1348gat));
  AOI21_X1  g733(.A(G176gat), .B1(new_n927), .B2(new_n615), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n930), .A2(new_n932), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n616), .B1(new_n372), .B2(new_n373), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1349gat));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n388), .A3(new_n675), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n930), .A2(new_n651), .A3(new_n932), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n358), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n356), .A3(new_n788), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n936), .A2(new_n636), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(G190gat), .ZN(new_n946));
  AOI211_X1 g745(.A(KEYINPUT61), .B(new_n356), .C1(new_n936), .C2(new_n636), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n530), .A2(new_n562), .A3(new_n549), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n925), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(KEYINPUT126), .B(G197gat), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n951), .A2(new_n729), .A3(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n932), .A2(new_n562), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n914), .B2(new_n915), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n862), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n949), .B(new_n955), .C1(new_n959), .C2(new_n952), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n952), .B1(new_n958), .B2(new_n862), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT127), .B1(new_n961), .B2(new_n954), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1352gat));
  NOR3_X1   g762(.A1(new_n951), .A2(G204gat), .A3(new_n616), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT62), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n616), .B(new_n957), .C1(new_n914), .C2(new_n915), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(new_n603), .ZN(G1353gat));
  INV_X1    g766(.A(new_n951), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n338), .A3(new_n675), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n958), .A2(new_n675), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AOI21_X1  g772(.A(G218gat), .B1(new_n968), .B2(new_n788), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n635), .A2(new_n339), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n958), .B2(new_n975), .ZN(G1355gat));
endmodule


