//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n470), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT65), .B1(new_n461), .B2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n461), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n468), .B1(new_n460), .B2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n476), .A2(new_n460), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT67), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n481), .A2(G124), .B1(G136), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n483), .A2(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(KEYINPUT68), .A2(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT68), .A2(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(G2104), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n476), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n463), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G102), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n471), .A2(new_n475), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n472), .A2(new_n474), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n460), .A2(G138), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT69), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n476), .B2(new_n498), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n465), .A2(new_n504), .A3(new_n499), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n514), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND2_X1  g097(.A1(new_n508), .A2(new_n510), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT70), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n527), .B1(new_n519), .B2(new_n528), .C1(new_n516), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n516), .A2(new_n534), .B1(new_n535), .B2(new_n519), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n533), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(new_n516), .ZN(new_n539));
  INV_X1    g114(.A(new_n519), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT71), .B(G43), .Z(new_n541));
  AOI22_X1  g116(.A1(new_n539), .A2(G81), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n513), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n540), .A2(KEYINPUT9), .A3(G53), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT9), .B1(new_n540), .B2(G53), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n539), .A2(G91), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n523), .B(KEYINPUT74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(KEYINPUT75), .B1(new_n564), .B2(G651), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n563), .A2(new_n566), .A3(new_n513), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n559), .B(new_n561), .C1(new_n565), .C2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n516), .A2(new_n571), .B1(new_n572), .B2(new_n519), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n511), .A2(G86), .A3(new_n515), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT76), .Z(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n523), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(G48), .A2(new_n540), .B1(new_n580), .B2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n516), .A2(new_n583), .B1(new_n584), .B2(new_n519), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n513), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n539), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  AOI22_X1  g166(.A1(new_n562), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n513), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n540), .A2(G54), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n589), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  XOR2_X1   g175(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g182(.A1(new_n481), .A2(G123), .B1(G135), .B2(new_n482), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G2096), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n465), .A2(new_n493), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XOR2_X1   g195(.A(G2427), .B(G2430), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G14), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(G401));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT18), .Z(new_n643));
  AOI21_X1  g218(.A(new_n639), .B1(KEYINPUT17), .B2(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n638), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n644), .B(new_n645), .C1(KEYINPUT17), .C2(new_n641), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n640), .B(KEYINPUT81), .Z(new_n647));
  OAI211_X1 g222(.A(new_n643), .B(new_n646), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(new_n612), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2100), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n661), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G1981), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  XOR2_X1   g246(.A(KEYINPUT82), .B(G29), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G35), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G162), .B2(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT93), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT29), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G19), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n546), .B2(new_n679), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n678), .A2(G2090), .B1(G1341), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n673), .A2(G26), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n481), .A2(G128), .B1(G140), .B2(new_n482), .ZN(new_n686));
  OR2_X1    g261(.A1(G104), .A2(G2105), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n687), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2067), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G16), .A2(G23), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT33), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G22), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G166), .B2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n697), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n697), .A2(KEYINPUT34), .A3(new_n702), .A4(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n482), .A2(G131), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT83), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n718), .A2(G95), .A3(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(G95), .B2(G2105), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n716), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n481), .B2(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(new_n673), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G25), .B2(new_n673), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT35), .B(G1991), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(G16), .A2(G24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G290), .B2(new_n679), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n711), .A2(new_n715), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n715), .B1(new_n711), .B2(new_n734), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n682), .B(new_n694), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n679), .A2(KEYINPUT23), .A3(G20), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n740));
  INV_X1    g315(.A(G20), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n742), .C1(new_n599), .C2(new_n679), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G1956), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G32), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT26), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n481), .B2(G129), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n493), .A2(G105), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G141), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(G29), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  AOI22_X1  g330(.A1(new_n744), .A2(new_n745), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n673), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n673), .ZN(new_n759));
  INV_X1    g334(.A(G2078), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n738), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n681), .A2(G1341), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n679), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n679), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n608), .A2(new_n610), .A3(new_n672), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G28), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n771), .A2(new_n772), .A3(new_n691), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n764), .A2(new_n768), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n679), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n679), .ZN(new_n777));
  INV_X1    g352(.A(G1961), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n679), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n595), .B2(new_n679), .ZN(new_n781));
  INV_X1    g356(.A(G1348), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n777), .A2(new_n778), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n779), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n744), .A2(new_n745), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n763), .A2(new_n775), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n493), .A2(G103), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT25), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n482), .A2(G139), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n793), .B(new_n794), .C1(new_n460), .C2(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G33), .B(new_n796), .S(G29), .Z(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT88), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  INV_X1    g374(.A(G2084), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G34), .ZN(new_n802));
  AOI22_X1  g377(.A1(G160), .A2(G29), .B1(new_n673), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n754), .A2(new_n755), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT91), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n678), .A2(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n800), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT92), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n790), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(G311));
  INV_X1    g386(.A(new_n790), .ZN(new_n812));
  INV_X1    g387(.A(new_n807), .ZN(new_n813));
  INV_X1    g388(.A(new_n808), .ZN(new_n814));
  INV_X1    g389(.A(new_n810), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(G150));
  NAND2_X1  g391(.A1(new_n540), .A2(G55), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n539), .A2(G93), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n817), .B(new_n818), .C1(new_n819), .C2(new_n513), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT95), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n595), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n546), .A2(new_n820), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT94), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n821), .A2(new_n544), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n546), .A2(new_n831), .A3(new_n820), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n827), .B(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n824), .B1(new_n834), .B2(G860), .ZN(G145));
  INV_X1    g410(.A(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n611), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(G162), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(G162), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n796), .A2(KEYINPUT97), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n752), .B(new_n723), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n690), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n482), .A2(G142), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT98), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n481), .A2(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n845), .A2(new_n690), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n846), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n853), .B1(new_n846), .B2(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n844), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n855), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n842), .B(new_n843), .C1(new_n859), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n503), .A2(new_n505), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n491), .A2(G2105), .B1(G102), .B2(new_n493), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n615), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n595), .B1(G299), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(G299), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n599), .A2(KEYINPUT99), .A3(new_n595), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n877), .A3(new_n873), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n833), .B(new_n604), .ZN(new_n880));
  MUX2_X1   g455(.A(new_n875), .B(new_n879), .S(new_n880), .Z(new_n881));
  XNOR2_X1  g456(.A(G305), .B(G288), .ZN(new_n882));
  XNOR2_X1  g457(.A(G290), .B(G303), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT101), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  MUX2_X1   g463(.A(new_n885), .B(new_n888), .S(KEYINPUT42), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n881), .B(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(KEYINPUT102), .A3(G868), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(G868), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(G868), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n822), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n892), .B2(new_n895), .ZN(G295));
  OAI21_X1  g471(.A(new_n891), .B1(new_n892), .B2(new_n895), .ZN(G331));
  NAND2_X1  g472(.A1(new_n833), .A2(G171), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n829), .A2(new_n830), .A3(G301), .A4(new_n832), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(G168), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G168), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n879), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n875), .A3(new_n900), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n884), .B(KEYINPUT100), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n867), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n903), .B2(new_n905), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n876), .A2(new_n912), .A3(new_n878), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n878), .A2(new_n912), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(new_n914), .C1(new_n901), .C2(new_n902), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n905), .ZN(new_n916));
  INV_X1    g491(.A(new_n906), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND4_X1   g493(.A1(KEYINPUT43), .A2(new_n918), .A3(new_n867), .A4(new_n907), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n918), .A2(new_n921), .A3(new_n867), .A4(new_n907), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n910), .B2(new_n921), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(G397));
  XNOR2_X1  g501(.A(KEYINPUT104), .B(G1384), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n864), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G160), .A2(G40), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n690), .B(G2067), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n752), .B(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n723), .B(new_n726), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(G290), .B2(G1986), .ZN(new_n940));
  OR3_X1    g515(.A1(G290), .A2(KEYINPUT105), .A3(G1986), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n932), .A2(G1986), .A3(G290), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT106), .Z(new_n945));
  NOR2_X1   g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G8), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n864), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n931), .B1(new_n949), .B2(new_n929), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n862), .B2(new_n863), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(KEYINPUT115), .A3(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT115), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n767), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(new_n931), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n951), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n800), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n947), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G168), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(new_n951), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(new_n947), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT109), .B(G1976), .Z(new_n969));
  NAND2_X1  g544(.A1(G288), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n699), .A2(G1976), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n967), .A2(new_n968), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(KEYINPUT110), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n577), .A2(new_n974), .A3(new_n581), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n581), .A2(new_n576), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G1981), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT49), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n967), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT111), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n967), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n968), .B1(new_n967), .B2(new_n971), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n972), .B1(new_n986), .B2(KEYINPUT110), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n973), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n950), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n705), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT107), .B(G2090), .Z(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n961), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n947), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G303), .A2(G8), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT55), .Z(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n964), .B1(new_n999), .B2(KEYINPUT116), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n995), .A2(new_n1003), .A3(new_n997), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n988), .B2(new_n998), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1000), .A2(KEYINPUT63), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n988), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n951), .A2(new_n959), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT112), .B1(new_n1011), .B2(new_n958), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n958), .B(KEYINPUT112), .C1(new_n951), .C2(new_n959), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT113), .B(new_n1010), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n993), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n960), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n957), .B1(new_n1018), .B2(new_n1013), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(KEYINPUT113), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n991), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n997), .B1(new_n1021), .B2(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1009), .B1(new_n1022), .B2(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g598(.A(new_n997), .ZN(new_n1024));
  INV_X1    g599(.A(new_n991), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n992), .B1(new_n1019), .B2(KEYINPUT113), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1010), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT114), .B(new_n1024), .C1(new_n1030), .C2(new_n947), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1023), .A2(new_n1032), .A3(new_n964), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1008), .B1(new_n1033), .B2(KEYINPUT63), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1005), .A2(new_n988), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n985), .A2(new_n1036), .A3(new_n699), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n975), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n967), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT126), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G168), .A2(new_n947), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n956), .B2(new_n962), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n952), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1966), .B1(new_n1048), .B2(new_n950), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1011), .A2(new_n958), .A3(new_n1010), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2084), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT121), .B(G8), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1043), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1043), .A2(KEYINPUT120), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1043), .A2(KEYINPUT120), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1052), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1044), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1041), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n955), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT122), .B(G1961), .Z(new_n1067));
  NAND2_X1  g642(.A1(new_n1050), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n950), .A2(new_n760), .A3(new_n989), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(KEYINPUT123), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT123), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1066), .B(new_n1068), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n963), .B2(KEYINPUT121), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(new_n1060), .B2(KEYINPUT51), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n1078), .C2(new_n1044), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1040), .A2(new_n1064), .A3(new_n1075), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1034), .A2(new_n1039), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n947), .B1(new_n1084), .B2(new_n991), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1083), .B1(new_n1085), .B2(new_n997), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(new_n1009), .A3(new_n1031), .A4(new_n1005), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1068), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(G301), .B(KEYINPUT54), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n930), .A2(new_n1092), .A3(new_n958), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(new_n989), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n930), .A2(new_n958), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1065), .B1(new_n1095), .B2(KEYINPUT124), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1090), .A2(new_n1097), .B1(new_n1073), .B2(new_n1091), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1078), .B2(new_n1044), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1082), .B1(new_n1087), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1027), .A2(new_n745), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n554), .A2(new_n556), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n561), .B(new_n1103), .C1(new_n565), .C2(new_n567), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n1105), .B2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(KEYINPUT117), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT57), .A3(G299), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n950), .A2(new_n989), .A3(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1101), .A2(new_n1106), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n966), .A2(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n965), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n990), .A2(G1996), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n546), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(G2067), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1115), .A2(new_n1122), .A3(new_n1117), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1050), .A2(new_n782), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n595), .ZN(new_n1129));
  INV_X1    g704(.A(new_n595), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1133), .A2(KEYINPUT60), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1113), .B(new_n1121), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1133), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1111), .A2(new_n595), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1108), .A2(new_n1106), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1073), .A2(new_n1091), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1097), .B(new_n1068), .C1(new_n1072), .C2(new_n1071), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1057), .A2(new_n1061), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1044), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1024), .B1(new_n1030), .B2(new_n947), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n988), .B1(new_n1148), .B2(new_n1083), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1031), .A2(new_n1005), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1147), .A2(KEYINPUT125), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1100), .A2(new_n1141), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n946), .B1(new_n1081), .B2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n942), .B(KEYINPUT48), .Z(new_n1154));
  NOR2_X1   g729(.A1(new_n939), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n937), .A2(new_n727), .A3(new_n723), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n690), .A2(new_n1122), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n933), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n753), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT127), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n935), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT46), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT47), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(KEYINPUT47), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1155), .B(new_n1158), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1153), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g742(.A(new_n650), .B1(new_n633), .B2(new_n634), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1169), .B1(new_n866), .B2(new_n867), .ZN(new_n1170));
  AND4_X1   g744(.A1(G319), .A2(new_n923), .A3(new_n1170), .A4(new_n670), .ZN(G308));
  NAND4_X1  g745(.A1(new_n923), .A2(new_n1170), .A3(G319), .A4(new_n670), .ZN(G225));
endmodule


