//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n461), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(new_n461), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n468), .A2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n475), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n475), .A2(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n461), .A2(KEYINPUT71), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n475), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n461), .A2(KEYINPUT71), .A3(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n460), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n491), .A2(new_n492), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  AND3_X1   g073(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT72), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n509), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n502), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n518), .A2(G651), .B1(G50), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n504), .A2(G89), .A3(new_n512), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n527), .B1(new_n499), .B2(new_n500), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT74), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n509), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n522), .A2(G51), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n526), .A2(new_n532), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  OAI211_X1 g113(.A(G52), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(G64), .B1(new_n499), .B2(new_n500), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n504), .A2(G90), .A3(new_n512), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(new_n513), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n516), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(G43), .B2(new_n522), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  AOI22_X1  g132(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G651), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n511), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n522), .A2(new_n564), .A3(G53), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n504), .A2(G91), .A3(new_n512), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n566), .A3(new_n567), .ZN(G299));
  NAND2_X1  g143(.A1(new_n544), .A2(new_n545), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n544), .A2(new_n545), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G301));
  NAND3_X1  g149(.A1(new_n504), .A2(G87), .A3(new_n512), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(KEYINPUT77), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(new_n580), .B1(G49), .B2(new_n522), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n577), .A2(KEYINPUT78), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT78), .B1(new_n577), .B2(new_n581), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n516), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n504), .A2(new_n512), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n522), .A2(G47), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n593), .B1(new_n559), .B2(new_n594), .C1(new_n591), .C2(new_n595), .ZN(G290));
  NAND3_X1  g171(.A1(new_n513), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n591), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  XOR2_X1   g176(.A(KEYINPUT80), .B(G66), .Z(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(new_n509), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n559), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n522), .A2(G54), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n607), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g183(.A(new_n607), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  NAND2_X1  g188(.A1(new_n604), .A2(new_n605), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(new_n597), .B2(new_n600), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n547), .A2(new_n551), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT81), .B1(new_n607), .B2(G559), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n615), .A2(new_n621), .A3(new_n616), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G868), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n481), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n483), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n461), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT84), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n460), .A2(new_n464), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n651), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n677), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(new_n674), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G33), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n460), .A2(G127), .ZN(new_n696));
  NAND2_X1  g271(.A1(G115), .A2(G2104), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n461), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n701));
  NAND3_X1  g276(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n481), .A2(G139), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n699), .A2(new_n700), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT99), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n695), .B1(new_n708), .B2(new_n694), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n709), .A2(G2072), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(G2072), .ZN(new_n711));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G5), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n569), .B2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G1961), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT102), .Z(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT30), .B(G28), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n718), .A2(new_n694), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n632), .B2(new_n694), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n712), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n712), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n722), .B1(G1966), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n717), .B(new_n725), .C1(G1966), .C2(new_n724), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n710), .B(new_n711), .C1(KEYINPUT103), .C2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n694), .A2(G32), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G129), .B2(new_n483), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT101), .Z(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G160), .B2(new_n694), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n694), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n694), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT106), .B(KEYINPUT29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2090), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G27), .A2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G164), .B2(G29), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT105), .B(G2078), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n737), .A2(new_n743), .A3(new_n748), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n694), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  AOI22_X1  g330(.A1(G128), .A2(new_n483), .B1(new_n481), .B2(G140), .ZN(new_n756));
  OAI21_X1  g331(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(G116), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n755), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT107), .B(KEYINPUT23), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n712), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1956), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n753), .A2(new_n764), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n712), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n552), .B2(new_n712), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n712), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n615), .B2(new_n712), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT93), .B(G1348), .Z(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n777), .A2(new_n779), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n774), .A2(new_n775), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n771), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  OAI22_X1  g358(.A1(new_n742), .A2(G2084), .B1(new_n734), .B2(new_n735), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n715), .B2(new_n714), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT104), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n726), .A2(KEYINPUT103), .ZN(new_n787));
  NOR4_X1   g362(.A1(new_n727), .A2(new_n783), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n712), .A2(G23), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n577), .A2(new_n581), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n791), .B2(new_n712), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT33), .B(G1976), .Z(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G6), .B(G305), .S(G16), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n712), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n712), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n792), .A2(new_n793), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n794), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n694), .A2(G25), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G131), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n483), .A2(G119), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n461), .A2(G107), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT89), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(G29), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT90), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n817), .ZN(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1986), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n805), .A2(new_n806), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  OR3_X1    g399(.A1(new_n823), .A2(KEYINPUT92), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n788), .A2(new_n825), .A3(new_n827), .ZN(G311));
  NAND3_X1  g403(.A1(new_n788), .A2(new_n825), .A3(new_n827), .ZN(G150));
  AOI22_X1  g404(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n559), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n504), .A2(G93), .A3(new_n512), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT109), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n522), .A2(G55), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n832), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n615), .A2(G559), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n552), .B(new_n831), .C1(new_n836), .C2(new_n835), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(new_n618), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n847), .B2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n839), .B1(new_n848), .B2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(new_n632), .B(new_n487), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G160), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n483), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n461), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(G142), .B2(new_n481), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n812), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n636), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n761), .B(new_n497), .ZN(new_n861));
  INV_X1    g436(.A(new_n733), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n707), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n707), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n863), .A2(new_n864), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n860), .B(new_n865), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  INV_X1    g447(.A(new_n860), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n870), .A3(new_n873), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n853), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n853), .A3(new_n869), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(G303), .B(KEYINPUT112), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n790), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT112), .ZN(new_n886));
  XNOR2_X1  g461(.A(G303), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n791), .ZN(new_n888));
  XNOR2_X1  g463(.A(G305), .B(G290), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n885), .B2(new_n888), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT42), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n615), .A2(new_n611), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n607), .A2(G299), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n843), .A2(new_n844), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n623), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n623), .A2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT111), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n894), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n615), .A2(new_n611), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n607), .A2(G299), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT41), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n900), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n898), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(new_n896), .C1(new_n899), .C2(new_n900), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n902), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT113), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n902), .A2(new_n915), .A3(new_n910), .A4(new_n912), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n893), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n893), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G868), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n837), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(G295));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n921), .ZN(G331));
  NAND3_X1  g498(.A1(new_n570), .A2(G168), .A3(new_n572), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n925));
  AND4_X1   g500(.A1(new_n925), .A2(G286), .A3(new_n545), .A4(new_n544), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(G171), .B2(G286), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT115), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n924), .B(KEYINPUT115), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n897), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT116), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT114), .B1(G168), .B2(new_n569), .ZN(new_n935));
  NAND3_X1  g510(.A1(G171), .A2(new_n925), .A3(G286), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT115), .B1(new_n937), .B2(new_n924), .ZN(new_n938));
  INV_X1    g513(.A(new_n931), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n845), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(KEYINPUT116), .A3(new_n897), .A4(new_n931), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n934), .A2(new_n896), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n932), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n897), .B1(new_n930), .B2(new_n931), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n908), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n892), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n879), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n890), .B2(new_n891), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT43), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n934), .A2(new_n940), .A3(new_n941), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n908), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n940), .A2(new_n896), .A3(new_n932), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n892), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n955), .A2(new_n947), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n956), .B1(new_n948), .B2(new_n950), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n955), .A2(new_n947), .A3(KEYINPUT43), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(KEYINPUT63), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n468), .A2(new_n479), .A3(G40), .ZN(new_n968));
  INV_X1    g543(.A(G2090), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n497), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n497), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n968), .A2(new_n969), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n468), .A2(new_n479), .A3(G40), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n975), .B1(new_n981), .B2(G1971), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n967), .B1(new_n982), .B2(G8), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n968), .A2(new_n977), .A3(new_n978), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n985), .A2(new_n975), .B1(new_n986), .B2(new_n800), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n972), .A2(new_n974), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n988), .A2(KEYINPUT118), .A3(new_n969), .A4(new_n968), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n990), .B2(new_n967), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n497), .A2(new_n970), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n992), .A2(G40), .A3(new_n468), .A4(new_n479), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT119), .A3(G8), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT119), .B1(new_n993), .B2(G8), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n790), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT120), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT120), .ZN(new_n1000));
  OAI221_X1 g575(.A(new_n1000), .B1(new_n997), .B2(new_n790), .C1(new_n995), .C2(new_n996), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(KEYINPUT52), .A3(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n582), .A2(new_n583), .A3(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT121), .B1(new_n1003), .B2(KEYINPUT52), .ZN(new_n1004));
  INV_X1    g579(.A(new_n998), .ZN(new_n1005));
  INV_X1    g580(.A(new_n583), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n577), .A2(KEYINPUT78), .A3(new_n581), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n997), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1005), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G305), .B(G1981), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(new_n996), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n994), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n991), .A2(new_n1002), .A3(new_n1012), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2084), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n988), .A2(new_n1019), .A3(new_n968), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n979), .B2(new_n980), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1023), .A2(G8), .A3(G168), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n964), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1002), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n987), .A2(new_n989), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n967), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n964), .B(new_n1024), .C1(new_n990), .C2(new_n967), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n560), .A2(new_n566), .A3(new_n567), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n979), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n968), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n972), .A2(new_n974), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n769), .B1(new_n1041), .B2(new_n980), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n968), .A2(new_n972), .A3(new_n974), .ZN(new_n1044));
  INV_X1    g619(.A(new_n993), .ZN(new_n1045));
  INV_X1    g620(.A(G2067), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(new_n778), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(new_n607), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1040), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n779), .B1(new_n988), .B2(new_n968), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n993), .A2(G2067), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n607), .B1(new_n1047), .B2(KEYINPUT60), .ZN(new_n1055));
  NOR4_X1   g630(.A1(new_n1052), .A2(new_n1053), .A3(new_n1051), .A4(new_n615), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1049), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1043), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT58), .B(G1341), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1045), .A2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT124), .B(G1996), .Z(new_n1063));
  NOR3_X1   g638(.A1(new_n979), .A2(new_n980), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n552), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT59), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n552), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1057), .A2(new_n1060), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1049), .B1(new_n1043), .B2(KEYINPUT125), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1040), .A2(new_n1037), .A3(new_n1072), .A4(new_n1042), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1050), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1002), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1076));
  INV_X1    g651(.A(new_n983), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1044), .A2(new_n715), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G2078), .ZN(new_n1082));
  OAI211_X1 g657(.A(G40), .B(new_n1082), .C1(new_n470), .C2(new_n461), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1083), .A2(new_n466), .A3(new_n467), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1038), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2078), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT53), .B1(new_n981), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(G171), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1081), .B1(new_n986), .B2(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n981), .A2(new_n1082), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(new_n1091), .A3(G301), .A4(new_n1080), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(KEYINPUT54), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT126), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT126), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1089), .A2(new_n1095), .A3(KEYINPUT54), .A4(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n1091), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n573), .B1(new_n1098), .B2(new_n1088), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(G301), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1086), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1023), .B2(G286), .ZN(new_n1103));
  AOI21_X1  g678(.A(G168), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(G8), .C1(new_n1023), .C2(G286), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1101), .A2(new_n1102), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1075), .A2(new_n1079), .A3(new_n1097), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(KEYINPUT62), .A3(new_n1107), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1099), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1079), .A3(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1017), .B(new_n997), .C1(new_n583), .C2(new_n582), .ZN(new_n1117));
  NOR2_X1   g692(.A1(G305), .A2(G1981), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT122), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n1016), .B1(new_n1026), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1033), .A2(new_n1109), .A3(new_n1116), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n980), .A2(new_n977), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(KEYINPUT117), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n761), .B(new_n1046), .ZN(new_n1126));
  INV_X1    g701(.A(G1996), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n733), .B(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n812), .B(new_n816), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G290), .B(G1986), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n813), .A2(new_n817), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(G2067), .B2(new_n761), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1125), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G290), .A2(G1986), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1125), .A2(KEYINPUT48), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1125), .A2(new_n1130), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT48), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT46), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT127), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1126), .A2(new_n862), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1144), .A2(new_n1145), .B1(new_n1125), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1150), .A2(KEYINPUT47), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT47), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1143), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1133), .A2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g729(.A1(new_n960), .A2(new_n961), .ZN(new_n1156));
  INV_X1    g730(.A(G319), .ZN(new_n1157));
  OR3_X1    g731(.A1(G401), .A2(G227), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g732(.A1(G229), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g733(.A(new_n1159), .B1(new_n877), .B2(new_n880), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1156), .A2(new_n1160), .ZN(G308));
  OAI221_X1 g735(.A(new_n1159), .B1(new_n877), .B2(new_n880), .C1(new_n960), .C2(new_n961), .ZN(G225));
endmodule


