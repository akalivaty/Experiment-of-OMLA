//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n212), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT67), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n212), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n228), .A2(G1), .A3(G13), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(new_n203), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n225), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n235), .B1(new_n220), .B2(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n222), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g0056(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n230), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n210), .A2(G33), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT11), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n209), .A2(G20), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G68), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n203), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT12), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(new_n265), .B2(KEYINPUT11), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G33), .A3(G41), .ZN(new_n281));
  INV_X1    g0081(.A(new_n226), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n284), .ZN(new_n288));
  INV_X1    g0088(.A(G238), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT76), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n228), .B1(G1), .B2(G13), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n278), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT70), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n227), .A2(new_n229), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(new_n278), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n239), .A2(G1698), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G226), .B2(G1698), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT3), .A2(G33), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n301), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n292), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n297), .B2(new_n278), .ZN(new_n309));
  AND2_X1   g0109(.A1(G33), .A2(G41), .ZN(new_n310));
  AOI211_X1 g0110(.A(KEYINPUT70), .B(new_n310), .C1(new_n227), .C2(new_n229), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n292), .B(new_n307), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n291), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT77), .A3(KEYINPUT13), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT77), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT76), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n290), .B1(new_n318), .B2(new_n312), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(new_n321), .A3(G179), .A4(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n322), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n323), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n327), .A2(new_n324), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n277), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n322), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n315), .A2(new_n321), .A3(G190), .A4(new_n322), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n332), .A2(new_n333), .A3(new_n276), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n337));
  INV_X1    g0137(.A(G226), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n287), .B1(new_n288), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT69), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT3), .B(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G222), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G223), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n344), .B1(new_n262), .B2(new_n342), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n300), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n339), .A2(new_n340), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n341), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT8), .B(G58), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT72), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(new_n263), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n356), .A2(new_n259), .B1(new_n201), .B2(new_n268), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n269), .A2(G50), .A3(new_n270), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT9), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n350), .A2(G200), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n357), .A2(KEYINPUT9), .A3(new_n358), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n352), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n350), .A2(new_n325), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(new_n359), .C1(G179), .C2(new_n350), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT73), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n354), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n263), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n259), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n269), .A2(G77), .A3(new_n270), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n268), .A2(new_n262), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n342), .A2(G232), .A3(new_n343), .ZN(new_n378));
  INV_X1    g0178(.A(G107), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n378), .B1(new_n379), .B2(new_n342), .C1(new_n345), .C2(new_n289), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n300), .ZN(new_n381));
  INV_X1    g0181(.A(new_n287), .ZN(new_n382));
  INV_X1    g0182(.A(new_n288), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n382), .B1(G244), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n377), .A2(KEYINPUT74), .B1(new_n385), .B2(G200), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n374), .A2(new_n375), .A3(new_n387), .A4(new_n376), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT75), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT75), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n391), .A3(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(new_n385), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G190), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G179), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n385), .A2(new_n325), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n377), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n338), .A2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G223), .B2(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G33), .ZN(new_n403));
  INV_X1    g0203(.A(G87), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n402), .A2(new_n306), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n300), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n382), .B1(G232), .B2(new_n383), .ZN(new_n407));
  AOI21_X1  g0207(.A(G169), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n396), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n306), .B2(new_n210), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  NOR4_X1   g0212(.A1(new_n304), .A2(new_n305), .A3(new_n412), .A4(G20), .ZN(new_n413));
  OAI21_X1  g0213(.A(G68), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(G58), .B(G68), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(KEYINPUT16), .A3(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n259), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n355), .B1(new_n209), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n269), .B1(new_n268), .B2(new_n355), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT18), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n410), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n406), .B2(new_n407), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n406), .A2(new_n407), .A3(G190), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n421), .A3(new_n423), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n430), .B1(G190), .B2(new_n409), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n421), .A4(new_n423), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n426), .A2(new_n428), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n400), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n337), .A2(new_n365), .A3(new_n369), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT82), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(G274), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n444), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n209), .A2(G45), .ZN(new_n452));
  INV_X1    g0252(.A(new_n448), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(new_n283), .A3(KEYINPUT82), .A4(G274), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n447), .B1(new_n449), .B2(new_n448), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n283), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n451), .A2(new_n456), .B1(new_n458), .B2(G257), .ZN(new_n459));
  OAI211_X1 g0259(.A(G244), .B(new_n343), .C1(new_n304), .C2(new_n305), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n342), .A2(KEYINPUT4), .A3(G244), .A4(new_n343), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n342), .A2(G250), .A3(G1698), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n300), .A2(new_n466), .A3(KEYINPUT81), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT81), .B1(new_n300), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n459), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n297), .B1(new_n256), .B2(new_n257), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n260), .A2(G77), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT6), .A2(G97), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(G97), .B(G107), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n472), .B1(new_n477), .B2(new_n210), .ZN(new_n478));
  OAI21_X1  g0278(.A(G107), .B1(new_n411), .B2(new_n413), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(KEYINPUT79), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n412), .B1(new_n342), .B2(G20), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n306), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n379), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n471), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n209), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n471), .A2(new_n487), .A3(new_n267), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n230), .A2(new_n258), .A3(new_n267), .A4(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT80), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n491), .A3(G97), .ZN(new_n492));
  INV_X1    g0292(.A(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n268), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n300), .A2(new_n466), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n459), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G190), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n470), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n206), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n503), .A2(KEYINPUT6), .B1(G107), .B2(new_n473), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n483), .B2(new_n484), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n259), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n494), .A3(new_n492), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n396), .B(new_n459), .C1(new_n467), .C2(new_n468), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n498), .A2(new_n325), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT83), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n452), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n209), .A2(new_n285), .A3(G45), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n513), .B1(new_n445), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n283), .A2(KEYINPUT83), .A3(new_n515), .A4(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n343), .C1(new_n304), .C2(new_n305), .ZN(new_n522));
  AND2_X1   g0322(.A1(KEYINPUT84), .A2(G116), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT84), .A2(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n521), .B(new_n522), .C1(new_n403), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n311), .B2(new_n309), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n520), .A2(new_n527), .A3(new_n396), .ZN(new_n528));
  AOI21_X1  g0328(.A(G169), .B1(new_n520), .B2(new_n527), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n372), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n489), .A2(new_n491), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n342), .A2(new_n210), .A3(G68), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n210), .B1(new_n301), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G87), .B2(new_n207), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n263), .B2(new_n493), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(new_n259), .B1(new_n268), .B2(new_n372), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n532), .A2(new_n533), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n533), .B1(new_n532), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n530), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n300), .A2(new_n526), .B1(new_n518), .B2(new_n519), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n520), .A2(new_n527), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n489), .A2(new_n491), .A3(G87), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n545), .A2(new_n547), .A3(new_n540), .A4(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n501), .A2(new_n512), .A3(new_n543), .A4(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n210), .B(G87), .C1(new_n304), .C2(new_n305), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT22), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT22), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n342), .A2(new_n553), .A3(new_n210), .A4(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n210), .B(G33), .C1(new_n523), .C2(new_n524), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT23), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n210), .B2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n379), .A2(KEYINPUT23), .A3(G20), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT86), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n555), .A2(KEYINPUT86), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(KEYINPUT24), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT86), .B1(new_n555), .B2(new_n561), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT24), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n471), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n489), .A2(new_n491), .A3(G107), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n268), .B(new_n379), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g0372(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n578));
  OAI211_X1 g0378(.A(G250), .B(new_n343), .C1(new_n304), .C2(new_n305), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G294), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n300), .A2(new_n581), .B1(G264), .B2(new_n458), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n451), .A2(new_n456), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n396), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n309), .B2(new_n311), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n458), .A2(G264), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n325), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT88), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n577), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n575), .B1(new_n566), .B2(new_n569), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n584), .A2(new_n588), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT88), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n587), .A2(new_n429), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n583), .A2(new_n585), .A3(new_n351), .A4(new_n586), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(new_n570), .A3(new_n576), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT89), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(KEYINPUT89), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n451), .A2(new_n456), .B1(new_n458), .B2(G270), .ZN(new_n605));
  OAI211_X1 g0405(.A(G264), .B(G1698), .C1(new_n304), .C2(new_n305), .ZN(new_n606));
  OAI211_X1 g0406(.A(G257), .B(new_n343), .C1(new_n304), .C2(new_n305), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n342), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n311), .B2(new_n309), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n325), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n471), .A2(G116), .A3(new_n267), .A4(new_n488), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n525), .A2(new_n268), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n403), .A2(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(G20), .B1(G33), .B2(G283), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n525), .A2(G20), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n259), .A2(KEYINPUT20), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT20), .B1(new_n259), .B2(new_n616), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n612), .B(new_n613), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(KEYINPUT21), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n619), .A2(G179), .A3(new_n610), .A4(new_n605), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT21), .B1(new_n611), .B2(new_n619), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n619), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n458), .A2(G270), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n610), .A2(new_n583), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G200), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n625), .B(new_n628), .C1(new_n351), .C2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NOR4_X1   g0430(.A1(new_n443), .A2(new_n550), .A3(new_n604), .A4(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n369), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n426), .A2(new_n428), .ZN(new_n633));
  INV_X1    g0433(.A(new_n330), .ZN(new_n634));
  INV_X1    g0434(.A(new_n399), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n335), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n437), .A2(new_n435), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n633), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n639), .B2(new_n365), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n543), .B(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n643));
  XNOR2_X1  g0443(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n543), .A3(new_n549), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n543), .A2(new_n549), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n646), .B2(new_n512), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n501), .A2(new_n512), .A3(new_n543), .A4(new_n549), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n577), .A2(new_n589), .A3(KEYINPUT90), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n592), .B2(new_n593), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n611), .A2(new_n619), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT21), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n621), .A3(new_n620), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n649), .B(new_n603), .C1(new_n653), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n640), .B1(new_n443), .B2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n625), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n630), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT93), .B(G330), .Z(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n577), .A2(new_n589), .A3(new_n667), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n592), .A2(new_n668), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n604), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n657), .A2(new_n668), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n595), .A3(new_n603), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n653), .A2(new_n668), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0486(.A(G41), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n223), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n233), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n659), .A2(new_n668), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n624), .A2(new_n591), .A3(new_n594), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n501), .A2(new_n512), .ZN(new_n697));
  INV_X1    g0497(.A(new_n646), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n603), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n543), .A4(new_n549), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n644), .B1(new_n646), .B2(new_n512), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n699), .A2(new_n642), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n695), .B1(new_n703), .B2(new_n668), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n544), .A2(new_n582), .A3(new_n459), .A4(new_n497), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n605), .A2(G179), .A3(new_n610), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n544), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n469), .A2(new_n587), .A3(new_n627), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(new_n711), .A3(KEYINPUT95), .ZN(new_n715));
  INV_X1    g0515(.A(new_n708), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n585), .A2(new_n586), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n546), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n499), .A3(new_n718), .A4(KEYINPUT30), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n714), .A2(new_n715), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n668), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n709), .A2(new_n711), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n667), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n720), .A2(new_n722), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n620), .A2(new_n621), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n656), .A3(new_n629), .A4(new_n668), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n649), .A2(new_n728), .A3(new_n595), .A4(new_n603), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n672), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n705), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n692), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(new_n688), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n210), .A2(G13), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n209), .B1(new_n736), .B2(G45), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n675), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n673), .B2(new_n671), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n223), .A2(new_n342), .ZN(new_n742));
  INV_X1    g0542(.A(G355), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n743), .B1(G116), .B2(new_n223), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n249), .A2(new_n446), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n223), .A2(new_n306), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n446), .B2(new_n234), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n744), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n230), .B1(G20), .B2(new_n325), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n210), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT96), .Z(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n739), .B1(new_n748), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT97), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n210), .A2(G190), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n210), .B1(new_n758), .B2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G97), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n396), .A2(G200), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G20), .A3(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n210), .A2(G179), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n429), .A2(G190), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n768), .A2(new_n202), .B1(new_n771), .B2(new_n379), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n351), .A2(new_n429), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n769), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(G87), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n210), .A2(new_n396), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n770), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n306), .B1(new_n779), .B2(G68), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n773), .A2(new_n777), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n759), .A2(new_n767), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(G50), .A2(new_n782), .B1(new_n784), .B2(G77), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n766), .A2(new_n776), .A3(new_n780), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n306), .B1(new_n774), .B2(new_n608), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT98), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n789), .B2(new_n760), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n765), .A2(G294), .ZN(new_n791));
  INV_X1    g0591(.A(new_n768), .ZN(new_n792));
  INV_X1    g0592(.A(new_n771), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G322), .B1(new_n793), .B2(G283), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n784), .A2(G311), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G326), .A2(new_n782), .B1(new_n779), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n791), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n763), .A2(new_n786), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n755), .B1(new_n799), .B2(new_n749), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n753), .B(KEYINPUT99), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n800), .B1(new_n671), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n741), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n751), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n750), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n739), .B1(new_n807), .B2(G77), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n768), .A2(new_n809), .B1(new_n783), .B2(new_n525), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n342), .B(new_n810), .C1(G107), .C2(new_n775), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n761), .A2(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n778), .A2(new_n813), .B1(new_n771), .B2(new_n404), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G303), .B2(new_n782), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n766), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n792), .A2(G143), .B1(new_n784), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n781), .C1(new_n819), .C2(new_n778), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT34), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n342), .B1(new_n771), .B2(new_n203), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n775), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n760), .B2(new_n824), .C1(new_n764), .C2(new_n202), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n816), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n808), .B1(new_n826), .B2(new_n749), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n399), .A2(new_n667), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n377), .A2(new_n667), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n395), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n399), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n827), .B1(new_n831), .B2(new_n806), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n395), .A2(new_n399), .A3(new_n668), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n657), .B1(new_n650), .B2(new_n652), .ZN(new_n834));
  AND4_X1   g0634(.A1(KEYINPUT89), .A2(new_n598), .A3(new_n570), .A4(new_n576), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT89), .B1(new_n592), .B2(new_n598), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n834), .A2(new_n837), .A3(new_n550), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT100), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n833), .B(new_n842), .C1(new_n838), .C2(new_n839), .ZN(new_n843));
  INV_X1    g0643(.A(new_n831), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n841), .A2(new_n843), .B1(new_n693), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n730), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n845), .A2(new_n730), .B1(new_n735), .B2(new_n738), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n832), .B1(new_n847), .B2(new_n848), .ZN(G384));
  OR2_X1    g0649(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(new_n851), .A3(G116), .A4(new_n231), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI211_X1 g0653(.A(new_n234), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n201), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n209), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n277), .A2(new_n667), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n330), .A2(new_n335), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n331), .A2(G169), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT14), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n327), .A2(new_n324), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n323), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n277), .B(new_n667), .C1(new_n863), .C2(new_n334), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n665), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n424), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n425), .A2(new_n433), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n665), .B1(new_n421), .B2(new_n423), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n870), .B2(KEYINPUT101), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n869), .B(new_n871), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n438), .A2(new_n870), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n869), .A2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n869), .A2(new_n871), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(KEYINPUT38), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n841), .A2(new_n843), .ZN(new_n880));
  INV_X1    g0680(.A(new_n828), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n866), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n872), .A2(new_n873), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n438), .A2(new_n870), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n869), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n877), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n330), .A2(new_n667), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n886), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n633), .A2(new_n867), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n442), .B1(new_n704), .B2(new_n694), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n640), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n898), .B(new_n900), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n724), .A2(KEYINPUT102), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT102), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n723), .A2(new_n903), .A3(new_n667), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(new_n721), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n723), .A2(new_n722), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n729), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT103), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n591), .A2(new_n594), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n837), .A2(new_n911), .A3(new_n727), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n649), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(KEYINPUT103), .A3(new_n905), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n844), .B1(new_n859), .B2(new_n864), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n891), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n865), .A2(new_n831), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n909), .B2(new_n914), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n879), .A2(KEYINPUT40), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n917), .A2(KEYINPUT40), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n442), .A2(new_n915), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n901), .B1(new_n672), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n209), .B2(new_n736), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n901), .A2(new_n672), .A3(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n857), .B1(new_n925), .B2(new_n926), .ZN(G367));
  INV_X1    g0727(.A(new_n754), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n223), .B2(new_n372), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n245), .A2(new_n746), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n739), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT109), .Z(new_n932));
  NAND3_X1  g0732(.A1(new_n775), .A2(KEYINPUT46), .A3(G116), .ZN(new_n933));
  INV_X1    g0733(.A(G311), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n933), .B1(new_n493), .B2(new_n771), .C1(new_n934), .C2(new_n781), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(G317), .B2(new_n761), .ZN(new_n936));
  INV_X1    g0736(.A(new_n525), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT46), .B1(new_n775), .B2(new_n937), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n608), .A2(new_n768), .B1(new_n778), .B2(new_n809), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n306), .B1(new_n783), .B2(new_n813), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n936), .B(new_n941), .C1(new_n379), .C2(new_n764), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT110), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n342), .B1(new_n771), .B2(new_n262), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT111), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n818), .B2(new_n760), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n764), .A2(new_n203), .ZN(new_n947));
  INV_X1    g0747(.A(G143), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n781), .A2(new_n948), .B1(new_n783), .B2(new_n201), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G150), .A2(new_n792), .B1(new_n779), .B2(G159), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n202), .B2(new_n774), .ZN(new_n951));
  NOR4_X1   g0751(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n943), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(KEYINPUT47), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n749), .B1(new_n953), .B2(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n548), .A2(new_n540), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n667), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n642), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT104), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n957), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n960), .B1(new_n646), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n958), .A2(new_n959), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n932), .B1(new_n954), .B2(new_n955), .C1(new_n964), .C2(new_n802), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n697), .B1(new_n496), .B2(new_n668), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n643), .A2(new_n667), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n679), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n682), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT42), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n911), .A2(new_n501), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n667), .B1(new_n975), .B2(new_n512), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n964), .A2(KEYINPUT105), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n962), .A2(KEYINPUT105), .A3(new_n963), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(KEYINPUT106), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT106), .B1(new_n982), .B2(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n982), .A2(new_n984), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT106), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(new_n970), .A3(new_n985), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n688), .B(KEYINPUT41), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n682), .B1(new_n678), .B2(new_n681), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n674), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n732), .A2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(KEYINPUT107), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n967), .A2(new_n968), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n684), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT44), .Z(new_n1002));
  INV_X1    g0802(.A(new_n679), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n684), .A2(new_n1000), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT45), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n998), .A2(new_n999), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n994), .B1(new_n1008), .B2(new_n733), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n993), .B(KEYINPUT108), .C1(new_n738), .C2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n992), .B(new_n988), .C1(new_n1009), .C2(new_n738), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT108), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n966), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n997), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(KEYINPUT114), .A3(new_n735), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n732), .A2(new_n996), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT114), .B1(new_n1016), .B2(new_n735), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n996), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n678), .A2(new_n802), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n742), .A2(new_n689), .B1(G107), .B2(new_n223), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n242), .A2(new_n446), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n689), .ZN(new_n1026));
  AOI211_X1 g0826(.A(G45), .B(new_n1026), .C1(G68), .C2(G77), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n354), .A2(G50), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n746), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1024), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n739), .B1(new_n1031), .B2(new_n754), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT112), .B(G150), .Z(new_n1033));
  INV_X1    g0833(.A(new_n355), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n761), .A2(new_n1033), .B1(new_n1034), .B2(new_n779), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n765), .A2(new_n531), .ZN(new_n1036));
  INV_X1    g0836(.A(G159), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1037), .A2(new_n781), .B1(new_n768), .B2(new_n201), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n774), .A2(new_n262), .B1(new_n783), .B2(new_n203), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n342), .B1(new_n771), .B2(new_n493), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1035), .A2(new_n1036), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G322), .A2(new_n782), .B1(new_n779), .B2(G311), .ZN(new_n1043));
  INV_X1    g0843(.A(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n608), .B2(new_n783), .C1(new_n1044), .C2(new_n768), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT113), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(KEYINPUT48), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n764), .A2(new_n813), .B1(new_n809), .B2(new_n774), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n306), .B1(new_n771), .B2(new_n525), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n761), .B2(G326), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1051), .A2(KEYINPUT49), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1042), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1032), .B1(new_n1057), .B2(new_n749), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1022), .A2(new_n738), .B1(new_n1023), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1021), .A2(new_n1059), .ZN(G393));
  AND2_X1   g0860(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1008), .B(new_n735), .C1(new_n997), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n738), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n928), .B1(new_n493), .B2(new_n223), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n252), .A2(new_n746), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n739), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n306), .B1(new_n771), .B2(new_n379), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G283), .A2(new_n775), .B1(new_n784), .B2(G294), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n608), .B2(new_n778), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G322), .C2(new_n761), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1044), .A2(new_n781), .B1(new_n768), .B2(new_n934), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n525), .C2(new_n764), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT115), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n765), .A2(G77), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n342), .B1(new_n771), .B2(new_n404), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n774), .A2(new_n203), .B1(new_n783), .B2(new_n354), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(G50), .C2(new_n779), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n761), .A2(G143), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n819), .A2(new_n781), .B1(new_n768), .B2(new_n1037), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1076), .A2(new_n1079), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1075), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1066), .B1(new_n1085), .B2(new_n749), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n753), .B2(new_n1000), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1062), .A2(new_n1063), .A3(new_n1087), .ZN(G390));
  NAND3_X1  g0888(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT39), .B1(new_n890), .B2(new_n877), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n879), .B2(KEYINPUT39), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n842), .B1(new_n659), .B2(new_n833), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n843), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n881), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n865), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n894), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1092), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n891), .A2(new_n1097), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n830), .A2(new_n399), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n703), .A2(new_n668), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n881), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1101), .B2(new_n881), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1099), .B1(new_n1105), .B2(new_n865), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1090), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n866), .B1(new_n731), .B2(new_n844), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1095), .ZN(new_n1110));
  AOI21_X1  g0910(.A(KEYINPUT103), .B1(new_n913), .B2(new_n905), .ZN(new_n1111));
  AND4_X1   g0911(.A1(KEYINPUT103), .A2(new_n905), .A3(new_n729), .A4(new_n906), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n831), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT117), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n866), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n730), .A2(new_n865), .A3(new_n831), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1101), .A2(new_n881), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1101), .A2(new_n1102), .A3(new_n881), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1114), .B1(new_n1113), .B2(new_n866), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1110), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n886), .A2(new_n893), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n866), .B1(new_n880), .B2(new_n881), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n894), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1118), .A2(new_n865), .A3(new_n1119), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1099), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n442), .A2(G330), .A3(new_n915), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n899), .A2(new_n1132), .A3(new_n640), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1107), .A2(new_n1123), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1113), .A2(new_n866), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT117), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1133), .B1(new_n1139), .B2(new_n1110), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT118), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1131), .A4(new_n1107), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1136), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1089), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1134), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n688), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1143), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1124), .A2(new_n751), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n739), .B1(new_n807), .B2(new_n1034), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT120), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n778), .A2(new_n379), .B1(new_n783), .B2(new_n493), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n761), .A2(G294), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n306), .B1(new_n774), .B2(new_n404), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n781), .A2(new_n813), .B1(new_n771), .B2(new_n203), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(G116), .C2(new_n792), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1154), .A2(new_n1153), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1076), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n342), .B1(new_n201), .B2(new_n771), .C1(new_n760), .C2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT119), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n775), .A2(new_n1033), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT53), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n765), .A2(G159), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G128), .A2(new_n782), .B1(new_n792), .B2(G132), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n779), .A2(G137), .B1(new_n784), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1160), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1152), .B1(new_n1172), .B2(new_n749), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1146), .A2(new_n738), .B1(new_n1151), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1150), .A2(new_n1174), .ZN(G378));
  NAND2_X1  g0975(.A1(new_n365), .A2(new_n367), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n359), .A2(new_n867), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n751), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n739), .B1(new_n807), .B2(G50), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n779), .A2(G97), .B1(new_n784), .B2(new_n531), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1184), .A2(KEYINPUT121), .B1(new_n760), .B2(new_n813), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n768), .A2(new_n379), .B1(new_n771), .B2(new_n202), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G116), .B2(new_n782), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G41), .B(new_n342), .C1(new_n775), .C2(G77), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n203), .C2(new_n764), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1185), .B(new_n1189), .C1(KEYINPUT121), .C2(new_n1184), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT122), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G33), .A2(G41), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1194), .C1(new_n306), .C2(new_n687), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n781), .A2(new_n1161), .B1(new_n778), .B2(new_n824), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G137), .B2(new_n784), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G128), .A2(new_n792), .B1(new_n775), .B2(new_n1169), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n819), .C2(new_n764), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  INV_X1    g1000(.A(G124), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1194), .B1(new_n1037), .B2(new_n771), .C1(new_n760), .C2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1199), .B2(KEYINPUT59), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1195), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1192), .A2(new_n1193), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1183), .B1(new_n1205), .B2(new_n749), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1182), .A2(new_n1206), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT123), .Z(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G330), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1181), .B1(new_n921), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n919), .A2(new_n920), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(G330), .A3(new_n1180), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1209), .B1(new_n1218), .B2(new_n737), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1135), .A2(KEYINPUT118), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1141), .B1(new_n1146), .B2(new_n1140), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1134), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1216), .B(new_n1217), .Z(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT57), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1133), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1125), .B1(new_n878), .B2(new_n874), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT125), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n896), .A4(new_n895), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1216), .A2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT125), .B1(new_n882), .B2(new_n897), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1215), .A3(new_n1211), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT57), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n735), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1220), .B1(new_n1225), .B2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1123), .A2(new_n738), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n739), .B1(new_n807), .B2(G68), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n774), .A2(new_n493), .B1(new_n783), .B2(new_n379), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n342), .B(new_n1240), .C1(G77), .C2(new_n793), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n761), .A2(G303), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n781), .A2(new_n809), .B1(new_n778), .B2(new_n525), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G283), .B2(new_n792), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1036), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n761), .A2(G128), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n768), .A2(new_n818), .B1(new_n783), .B2(new_n819), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G132), .B2(new_n782), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n306), .B1(new_n793), .B2(G58), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G159), .A2(new_n775), .B1(new_n779), .B2(new_n1169), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n764), .A2(new_n201), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1239), .B1(new_n1253), .B2(new_n749), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n865), .B2(new_n806), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1238), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n994), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1139), .A2(new_n1110), .A3(new_n1133), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1148), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(G381));
  INV_X1    g1061(.A(G381), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n804), .B(new_n1059), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(G390), .A2(G384), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1014), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT57), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1226), .B2(new_n1218), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1223), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1269), .A3(new_n735), .ZN(new_n1270));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1220), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1265), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1273), .B(new_n1274), .ZN(G407));
  NOR2_X1   g1075(.A1(new_n1272), .A2(G343), .ZN(new_n1276));
  INV_X1    g1076(.A(G213), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G407), .A2(new_n1278), .ZN(G409));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1280), .A2(G390), .A3(new_n1263), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1063), .A2(new_n1087), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n804), .B1(new_n1021), .B2(new_n1059), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1263), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1062), .B(new_n1282), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1014), .B(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G375), .A2(G378), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT62), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1291), .A2(new_n1259), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1139), .A2(KEYINPUT60), .A3(new_n1110), .A4(new_n1133), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n735), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G384), .B(new_n1257), .C1(new_n1292), .C2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(G384), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1291), .B2(new_n1259), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1256), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1207), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1234), .B2(new_n738), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1150), .A2(new_n1302), .A3(new_n1174), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1223), .A2(new_n1258), .A3(new_n1224), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n1303), .A2(new_n1304), .B1(G213), .B2(new_n666), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1289), .A2(new_n1290), .A3(new_n1300), .A4(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1295), .A2(new_n1298), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1271), .B1(new_n1270), .B2(new_n1220), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1150), .A2(new_n1302), .A3(new_n1174), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1226), .A2(new_n1218), .A3(new_n994), .ZN(new_n1313));
  OAI22_X1  g1113(.A1(new_n1312), .A2(new_n1313), .B1(new_n1277), .B2(G343), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1310), .B1(new_n1311), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1306), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1314), .B1(G378), .B2(G375), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(new_n1300), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1288), .B1(new_n1317), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1289), .A2(new_n1305), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1323), .B2(new_n1299), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1310), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1287), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1321), .A2(new_n1327), .ZN(G405));
  NAND2_X1  g1128(.A1(new_n1289), .A2(new_n1272), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1300), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1289), .A2(new_n1272), .A3(new_n1299), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1287), .A2(new_n1330), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1287), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(G402));
endmodule


