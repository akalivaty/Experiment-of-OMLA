//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT0), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n206), .A2(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G68), .A2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(KEYINPUT64), .A2(G77), .ZN(new_n222));
  NOR2_X1   g0022(.A1(KEYINPUT64), .A2(G77), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n221), .B1(G244), .B2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n229), .B(new_n230), .C1(new_n226), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n207), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n216), .B1(new_n206), .B2(new_n209), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n255), .A2(new_n252), .A3(G13), .A4(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n213), .B1(new_n207), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT69), .Z(new_n262));
  AOI21_X1  g0062(.A(new_n202), .B1(new_n252), .B2(G20), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n214), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n257), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n270), .A2(new_n259), .B1(new_n202), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n282), .B2(G226), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(G223), .A3(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G222), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n289), .B1(new_n224), .B2(new_n288), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n275), .B(new_n296), .C1(new_n297), .C2(new_n295), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n274), .A2(KEYINPUT9), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n295), .A2(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(G200), .B2(new_n295), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n299), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n275), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n295), .A2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n273), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n288), .A2(G232), .A3(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(new_n291), .C2(new_n218), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n279), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n278), .B1(new_n282), .B2(G238), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n312), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n320), .A2(G190), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n318), .B2(KEYINPUT73), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  AOI211_X1 g0125(.A(new_n325), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n326));
  OAI21_X1  g0126(.A(G200), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n261), .B1(new_n252), .B2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G68), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT75), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n271), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT12), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n266), .A2(G50), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(new_n214), .B2(G68), .ZN(new_n335));
  INV_X1    g0135(.A(G77), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n269), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n259), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT11), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n323), .A2(new_n327), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G169), .B1(new_n324), .B2(new_n326), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(G169), .C1(new_n324), .C2(new_n326), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n320), .A2(G179), .A3(new_n321), .A4(new_n322), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n341), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n328), .A2(G77), .ZN(new_n353));
  INV_X1    g0153(.A(new_n266), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n224), .A2(new_n214), .B1(new_n268), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n269), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n259), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n271), .A2(new_n224), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n288), .A2(G238), .A3(G1698), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n288), .A2(G232), .A3(new_n290), .ZN(new_n362));
  INV_X1    g0162(.A(G107), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n288), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n279), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n278), .B1(new_n282), .B2(G244), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(new_n369), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n360), .B1(new_n371), .B2(G169), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n308), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n372), .A2(new_n373), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n360), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n371), .A2(G200), .ZN(new_n380));
  AOI21_X1  g0180(.A(G190), .B1(new_n368), .B2(new_n370), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n311), .A2(new_n352), .A3(new_n378), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT84), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n281), .A2(new_n386), .B1(new_n277), .B2(new_n276), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT76), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n258), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT76), .A2(G33), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(KEYINPUT3), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n286), .ZN(new_n393));
  NAND2_X1  g0193(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(G33), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n290), .A2(G223), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n218), .B2(new_n290), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n387), .B1(new_n401), .B2(new_n279), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n308), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G169), .B2(new_n402), .ZN(new_n404));
  XOR2_X1   g0204(.A(new_n404), .B(KEYINPUT82), .Z(new_n405));
  INV_X1    g0205(.A(KEYINPUT81), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT78), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n391), .A2(new_n395), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n214), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G68), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n409), .B1(new_n408), .B2(new_n214), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT7), .B1(new_n396), .B2(G20), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT78), .A3(G68), .A4(new_n410), .ZN(new_n415));
  XNOR2_X1  g0215(.A(G58), .B(G68), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(G20), .B1(G159), .B2(new_n266), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT16), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n259), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT80), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n421));
  AND2_X1   g0221(.A1(KEYINPUT76), .A2(G33), .ZN(new_n422));
  NOR2_X1   g0222(.A1(KEYINPUT76), .A2(G33), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n286), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(KEYINPUT79), .B1(new_n425), .B2(new_n258), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n286), .C1(new_n422), .C2(new_n423), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n285), .A2(new_n287), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT7), .B1(new_n430), .B2(new_n214), .ZN(new_n431));
  OAI21_X1  g0231(.A(G68), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n420), .B(KEYINPUT16), .C1(new_n432), .C2(new_n417), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n424), .A2(KEYINPUT79), .ZN(new_n434));
  INV_X1    g0234(.A(new_n394), .ZN(new_n435));
  NOR2_X1   g0235(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n258), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n421), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n417), .B1(new_n440), .B2(new_n331), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT16), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT80), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n419), .A2(new_n433), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n268), .B1(new_n252), .B2(G20), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n262), .A2(new_n445), .B1(new_n271), .B2(new_n268), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n406), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT3), .B1(new_n389), .B2(new_n390), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n437), .B1(new_n449), .B2(new_n427), .ZN(new_n450));
  INV_X1    g0250(.A(new_n428), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n431), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n331), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n417), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n442), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n420), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n441), .A2(KEYINPUT80), .A3(new_n442), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n457), .A2(new_n259), .A3(new_n418), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT81), .A3(new_n446), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n405), .A2(new_n448), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n405), .A2(new_n448), .A3(KEYINPUT18), .A4(new_n460), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n402), .A2(new_n297), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G200), .B2(new_n402), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n459), .A2(new_n446), .A3(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n467), .A2(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT83), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n459), .A2(new_n470), .A3(new_n446), .A4(new_n466), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(KEYINPUT17), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n463), .A2(new_n464), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n384), .A2(new_n385), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n385), .B1(new_n384), .B2(new_n473), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G264), .A2(G1698), .ZN(new_n478));
  OR3_X1    g0278(.A1(new_n408), .A2(KEYINPUT87), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n430), .A2(G303), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n396), .A2(G257), .A3(new_n290), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT87), .B1(new_n408), .B2(new_n478), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n279), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT88), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n279), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G41), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n252), .B(G45), .C1(new_n489), .C2(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT85), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(KEYINPUT5), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(G274), .A3(new_n280), .A4(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n493), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n490), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n279), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(G270), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n261), .B1(new_n252), .B2(G33), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  INV_X1    g0303(.A(G97), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n504), .B2(G33), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n214), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G20), .A2(G116), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n260), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n271), .A2(new_n219), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G169), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n500), .A2(new_n513), .A3(KEYINPUT21), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  INV_X1    g0315(.A(new_n499), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n486), .B2(new_n487), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(G179), .A3(new_n511), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G200), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n500), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n297), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n511), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  MUX2_X1   g0325(.A(G250), .B(G257), .S(G1698), .Z(new_n526));
  NAND2_X1  g0326(.A1(new_n396), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n389), .A2(new_n390), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G294), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n280), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n498), .A2(G264), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n495), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G179), .ZN(new_n534));
  INV_X1    g0334(.A(G169), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n533), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT89), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  INV_X1    g0338(.A(G87), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n396), .A2(new_n214), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n214), .A2(G87), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n430), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n528), .A2(new_n214), .A3(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n214), .A2(G107), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT23), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n547), .B2(KEYINPUT24), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(KEYINPUT24), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n547), .A2(new_n537), .A3(KEYINPUT24), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n260), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n501), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT25), .B1(new_n257), .B2(G107), .ZN(new_n555));
  OR3_X1    g0355(.A1(new_n257), .A2(KEYINPUT25), .A3(G107), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n536), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n530), .A2(new_n532), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n297), .A3(new_n494), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G200), .B2(new_n533), .ZN(new_n561));
  INV_X1    g0361(.A(new_n557), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n551), .A2(new_n548), .A3(new_n549), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n260), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT90), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n558), .A2(KEYINPUT90), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(G107), .B1(new_n429), .B2(new_n431), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n363), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n504), .A2(new_n363), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n571), .B1(new_n574), .B2(KEYINPUT6), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n260), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n257), .A2(G97), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n501), .B2(G97), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n396), .A2(G244), .A3(new_n290), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT4), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n288), .A2(G250), .A3(G1698), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n585), .A2(new_n503), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n280), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n498), .A2(G257), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n494), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n588), .A2(G190), .A3(new_n590), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n581), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G169), .B1(new_n588), .B2(new_n590), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n494), .A2(new_n589), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n503), .A3(new_n586), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n583), .B2(new_n582), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(G179), .C1(new_n598), .C2(new_n280), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n577), .B2(new_n580), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n396), .A2(new_n214), .A3(G68), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n214), .B1(new_n314), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G87), .A2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n363), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n606), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n260), .B1(new_n602), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n356), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n257), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n501), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n396), .A2(G238), .A3(new_n290), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n396), .A2(G244), .A3(G1698), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n528), .A2(G116), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n279), .ZN(new_n619));
  INV_X1    g0419(.A(G45), .ZN(new_n620));
  OAI21_X1  g0420(.A(G250), .B1(new_n620), .B2(G1), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n252), .A2(G45), .A3(G274), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n279), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n619), .A2(new_n308), .A3(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n618), .A2(new_n279), .B1(new_n624), .B2(new_n625), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n614), .B(new_n627), .C1(G169), .C2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n619), .A2(G190), .A3(new_n626), .ZN(new_n630));
  AOI211_X1 g0430(.A(new_n539), .B(new_n261), .C1(new_n252), .C2(G33), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n631), .A2(new_n609), .A3(new_n611), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(new_n632), .C1(new_n521), .C2(new_n628), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n594), .A2(new_n601), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n477), .A2(new_n525), .A3(new_n569), .A4(new_n634), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n472), .A2(new_n468), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n349), .A2(new_n350), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n636), .B(new_n342), .C1(new_n638), .C2(new_n378), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n404), .B1(new_n459), .B2(new_n446), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n306), .B1(new_n273), .B2(new_n309), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n634), .A2(new_n564), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n558), .A2(new_n514), .A3(new_n518), .A4(new_n519), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n629), .A2(new_n633), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n581), .B1(new_n599), .B2(new_n595), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g0450(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n651));
  OAI21_X1  g0451(.A(new_n629), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n643), .B1(new_n476), .B2(new_n656), .ZN(G369));
  NAND3_X1  g0457(.A1(new_n252), .A2(new_n214), .A3(G13), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n553), .B2(new_n557), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n569), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n663), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n558), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n511), .A2(new_n663), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n520), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n520), .B2(new_n524), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n520), .A2(new_n666), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n665), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n558), .A2(new_n663), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n208), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n605), .A2(new_n363), .A3(new_n219), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n211), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT28), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT93), .B1(new_n656), .B2(new_n663), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n663), .B1(new_n646), .B2(new_n655), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AND4_X1   g0494(.A1(new_n564), .A2(new_n594), .A3(new_n601), .A4(new_n633), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n645), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n651), .B1(new_n647), .B2(new_n601), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n649), .A2(new_n653), .A3(new_n629), .A4(new_n633), .ZN(new_n698));
  AND3_X1   g0498(.A1(new_n697), .A2(new_n629), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n663), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n569), .A2(new_n525), .A3(new_n634), .A4(new_n666), .ZN(new_n703));
  NOR4_X1   g0503(.A1(new_n591), .A2(new_n533), .A3(new_n628), .A4(G179), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n500), .ZN(new_n705));
  XOR2_X1   g0505(.A(new_n705), .B(KEYINPUT92), .Z(new_n706));
  AND3_X1   g0506(.A1(new_n591), .A2(new_n559), .A3(new_n628), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n517), .A2(new_n707), .A3(G179), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n703), .A2(KEYINPUT31), .B1(new_n710), .B2(new_n663), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  AOI211_X1 g0512(.A(new_n712), .B(new_n666), .C1(new_n709), .C2(new_n705), .ZN(new_n713));
  OAI21_X1  g0513(.A(G330), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n702), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n688), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(G13), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n685), .B1(G45), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n674), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n672), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n521), .A2(G179), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G20), .A3(G190), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G87), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n214), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n730), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n288), .C1(new_n363), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT96), .Z(new_n737));
  NAND2_X1  g0537(.A1(G20), .A2(G179), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT95), .Z(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n297), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n521), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(G200), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n737), .B1(new_n331), .B2(new_n742), .C1(new_n224), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n297), .A2(new_n521), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G50), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n297), .A2(G200), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n739), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G58), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n734), .A2(new_n754), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n749), .A2(new_n753), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n742), .A2(new_n763), .B1(new_n751), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  INV_X1    g0566(.A(G326), .ZN(new_n767));
  INV_X1    g0567(.A(new_n756), .ZN(new_n768));
  INV_X1    g0568(.A(G294), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n747), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n743), .A2(G311), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n731), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n430), .B1(new_n735), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n758), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n775), .B(new_n777), .C1(G329), .C2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n745), .A2(new_n762), .B1(new_n766), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n213), .B1(G20), .B2(new_n535), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n288), .A2(G355), .A3(new_n208), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G116), .B2(new_n208), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n247), .A2(G45), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n212), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n396), .A2(new_n682), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n727), .A2(new_n782), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n720), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT94), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n783), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n722), .A2(new_n724), .B1(new_n729), .B2(new_n794), .ZN(G396));
  NOR2_X1   g0595(.A1(new_n782), .A2(new_n725), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n219), .A2(new_n744), .B1(new_n742), .B2(new_n776), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n769), .A2(new_n751), .B1(new_n747), .B2(new_n774), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n288), .B1(new_n778), .B2(G311), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n732), .A2(G107), .ZN(new_n801));
  INV_X1    g0601(.A(new_n735), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G87), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n800), .A2(new_n801), .A3(new_n757), .A4(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n798), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G137), .A2(new_n748), .B1(new_n752), .B2(G143), .ZN(new_n806));
  INV_X1    g0606(.A(G150), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n742), .B2(new_n807), .C1(new_n759), .C2(new_n744), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(G68), .ZN(new_n810));
  INV_X1    g0610(.A(G132), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n202), .B2(new_n731), .C1(new_n811), .C2(new_n758), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n408), .B(new_n812), .C1(G58), .C2(new_n756), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n805), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n782), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n720), .B1(G77), .B2(new_n797), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT99), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n360), .A2(new_n663), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n376), .A2(new_n377), .B1(new_n382), .B2(new_n818), .ZN(new_n819));
  AND4_X1   g0619(.A1(new_n377), .A2(new_n374), .A3(new_n375), .A4(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n817), .B1(new_n726), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n690), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n689), .A2(new_n692), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n821), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n825), .A2(new_n714), .ZN(new_n826));
  INV_X1    g0626(.A(new_n720), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n825), .B2(new_n714), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n826), .B2(new_n828), .ZN(G384));
  AOI21_X1  g0629(.A(new_n224), .B1(G58), .B2(G68), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(new_n212), .B1(new_n202), .B2(G68), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n831), .A2(new_n252), .A3(G13), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT101), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n215), .A2(G116), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n575), .B(KEYINPUT100), .Z(new_n835));
  INV_X1    g0635(.A(KEYINPUT35), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT36), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n712), .B(new_n666), .C1(new_n706), .C2(new_n709), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n711), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n350), .A2(new_n663), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n637), .A2(KEYINPUT102), .A3(new_n342), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n349), .A2(new_n350), .A3(new_n663), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT102), .B1(new_n351), .B2(new_n844), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n843), .A2(new_n821), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT104), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n459), .A2(new_n446), .A3(new_n466), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n640), .ZN(new_n856));
  INV_X1    g0656(.A(new_n661), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n448), .A2(new_n460), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n433), .A2(new_n443), .ZN(new_n859));
  INV_X1    g0659(.A(new_n419), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n447), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n467), .B(KEYINPUT104), .C1(new_n861), .C2(new_n404), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n856), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n469), .A2(new_n865), .A3(new_n471), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n448), .B(new_n460), .C1(new_n405), .C2(new_n857), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n864), .A2(KEYINPUT105), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n636), .A2(new_n641), .ZN(new_n870));
  INV_X1    g0670(.A(new_n858), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n863), .A2(KEYINPUT37), .B1(new_n866), .B2(new_n867), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n853), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n415), .A2(new_n417), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT16), .B1(new_n877), .B2(new_n413), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n446), .B1(new_n878), .B2(new_n419), .ZN(new_n879));
  INV_X1    g0679(.A(new_n404), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n879), .B1(new_n880), .B2(new_n857), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n469), .A2(new_n471), .A3(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n866), .A2(new_n867), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n857), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n884), .B(KEYINPUT38), .C1(new_n473), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n852), .A2(KEYINPUT40), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n463), .A2(new_n464), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n889), .B2(new_n636), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n853), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n886), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT40), .B1(new_n852), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n477), .A2(new_n843), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n894), .B(new_n895), .Z(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(G330), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT106), .Z(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n891), .B2(new_n886), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n890), .A2(new_n853), .A3(new_n883), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n858), .B1(new_n636), .B2(new_n641), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n874), .B2(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n864), .A2(new_n868), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n901), .B1(new_n907), .B2(new_n853), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n900), .B1(new_n908), .B2(new_n899), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n637), .A2(new_n663), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n376), .A2(new_n377), .A3(new_n666), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n690), .B2(new_n821), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n892), .A2(new_n916), .A3(new_n850), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n641), .B2(new_n857), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n694), .B(new_n701), .C1(new_n474), .C2(new_n475), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n643), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n898), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(G1), .B1(new_n718), .B2(G20), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n898), .B2(new_n922), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT107), .B1(new_n923), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n841), .B1(new_n926), .B2(new_n927), .ZN(G367));
  INV_X1    g0728(.A(new_n788), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n243), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n791), .B1(new_n682), .B2(new_n610), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n827), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n756), .A2(G68), .ZN(new_n934));
  AOI22_X1  g0734(.A1(G143), .A2(new_n748), .B1(new_n752), .B2(G150), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n430), .B1(new_n732), .B2(G58), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n225), .A2(new_n802), .B1(new_n778), .B2(G137), .ZN(new_n937));
  AND4_X1   g0737(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n202), .B2(new_n744), .C1(new_n759), .C2(new_n742), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n802), .A2(G97), .B1(new_n778), .B2(G317), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n408), .C1(new_n774), .C2(new_n751), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(G311), .B2(new_n748), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n732), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT46), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n731), .B2(new_n219), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n945), .C1(new_n363), .C2(new_n768), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n741), .B2(G294), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n942), .B(new_n947), .C1(new_n776), .C2(new_n744), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n939), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT47), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n782), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(KEYINPUT47), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n632), .A2(new_n666), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n648), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n629), .B2(new_n953), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n933), .B1(new_n951), .B2(new_n952), .C1(new_n728), .C2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n667), .A2(new_n674), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n677), .B1(new_n675), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n665), .A2(new_n677), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n702), .A2(new_n959), .A3(new_n714), .A4(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n960), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n965), .A2(KEYINPUT111), .A3(new_n714), .A4(new_n702), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n594), .B(new_n601), .C1(new_n581), .C2(new_n666), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n649), .A2(new_n663), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT44), .B1(new_n680), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  INV_X1    g0772(.A(new_n970), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(new_n678), .C2(new_n679), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n680), .B2(new_n970), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n971), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n676), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(KEYINPUT110), .A3(new_n675), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n716), .B1(new_n967), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT112), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n683), .B(KEYINPUT41), .Z(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n977), .A2(KEYINPUT110), .A3(new_n675), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n675), .B1(new_n977), .B2(KEYINPUT110), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n963), .A2(new_n966), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n715), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT112), .B1(new_n991), .B2(new_n984), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n719), .A2(G45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(G1), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n986), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n960), .A2(new_n968), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n601), .B1(new_n968), .B2(new_n558), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n997), .A2(KEYINPUT42), .B1(new_n666), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n955), .B(KEYINPUT43), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT109), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n999), .A2(new_n1007), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1009), .A2(new_n1011), .B1(new_n676), .B2(new_n973), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1008), .A2(new_n1006), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n676), .A2(new_n973), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1013), .A2(new_n1014), .A3(new_n1010), .A4(new_n1005), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n957), .B1(new_n996), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(G387));
  NAND2_X1  g0818(.A1(new_n715), .A2(new_n964), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n683), .A3(new_n961), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n331), .A2(new_n744), .B1(new_n742), .B2(new_n268), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n732), .A2(new_n225), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n802), .A2(G97), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n778), .A2(G150), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n396), .A4(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT114), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n768), .A2(new_n356), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n752), .B2(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n759), .B2(new_n747), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1021), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n735), .A2(new_n219), .B1(new_n758), .B2(new_n767), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n752), .B1(new_n748), .B2(G322), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n774), .B2(new_n744), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G311), .B2(new_n741), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT48), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(KEYINPUT48), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n732), .A2(G294), .B1(new_n756), .B2(G283), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n396), .B(new_n1031), .C1(new_n1039), .C2(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(KEYINPUT49), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n815), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n667), .A2(new_n728), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n268), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n686), .C1(G68), .C2(G77), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n929), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n239), .B2(new_n620), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n288), .A2(new_n208), .A3(new_n686), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(G107), .B2(new_n208), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT113), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n791), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1043), .A2(new_n1044), .A3(new_n827), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n965), .B2(new_n994), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1020), .A2(new_n1055), .ZN(G393));
  OR2_X1    g0856(.A1(new_n977), .A2(new_n676), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n977), .A2(new_n676), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n961), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n683), .C1(new_n967), .C2(new_n981), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n994), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n790), .B1(new_n504), .B2(new_n208), .C1(new_n929), .C2(new_n250), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n720), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n752), .B1(new_n748), .B2(G317), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n430), .B1(new_n735), .B2(new_n363), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n731), .A2(new_n776), .B1(new_n758), .B2(new_n764), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G116), .C2(new_n756), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n742), .B2(new_n774), .C1(new_n769), .C2(new_n744), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n803), .B1(new_n331), .B2(new_n731), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n768), .A2(new_n336), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n778), .A2(G143), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .A4(new_n408), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n202), .B2(new_n742), .C1(new_n268), .C2(new_n744), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n807), .A2(new_n747), .B1(new_n751), .B2(new_n759), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT51), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n1066), .A2(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1064), .B1(new_n1078), .B2(new_n782), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n970), .B2(new_n728), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1060), .A2(new_n1062), .A3(new_n1080), .ZN(G390));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n914), .B1(new_n700), .B2(new_n821), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n912), .B1(new_n1083), .B2(new_n849), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n908), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1084), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n887), .A2(KEYINPUT115), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n876), .A2(new_n899), .A3(new_n886), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n900), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n912), .B1(new_n915), .B2(new_n849), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  OAI211_X1 g0892(.A(G330), .B(new_n821), .C1(new_n711), .C2(new_n713), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n850), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1088), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1085), .A2(new_n1087), .B1(new_n909), .B2(new_n1091), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n821), .C1(new_n711), .C2(new_n842), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n849), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(KEYINPUT116), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT115), .B1(new_n887), .B2(new_n1086), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1082), .B(new_n1084), .C1(new_n876), .C2(new_n886), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1092), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT116), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n1100), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1097), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n994), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n909), .A2(new_n725), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n827), .B1(new_n268), .B2(new_n796), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n741), .A2(G137), .B1(G159), .B2(new_n756), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1112), .B1(new_n744), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT119), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n732), .A2(G150), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1118), .A2(new_n747), .B1(new_n751), .B2(new_n811), .ZN(new_n1119));
  INV_X1    g0919(.A(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n288), .B1(new_n758), .B2(new_n1120), .C1(new_n202), .C2(new_n735), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n219), .A2(new_n751), .B1(new_n747), .B2(new_n776), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n778), .A2(G294), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n733), .A2(new_n810), .A3(new_n1124), .A4(new_n430), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1123), .A2(new_n1125), .A3(new_n1072), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G97), .A2(new_n743), .B1(new_n741), .B2(G107), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1115), .A2(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1110), .B(new_n1111), .C1(new_n815), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1109), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n843), .B(G330), .C1(new_n474), .C2(new_n475), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n920), .A2(new_n1131), .A3(new_n643), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1099), .A2(new_n849), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1083), .B1(new_n1093), .B2(new_n849), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT117), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT117), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1095), .A2(new_n1137), .A3(new_n1083), .A4(new_n1133), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1094), .A2(new_n850), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n916), .B1(new_n1140), .B2(new_n1100), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1132), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1108), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n684), .ZN(new_n1144));
  AOI211_X1 g0944(.A(KEYINPUT116), .B(new_n1101), .C1(new_n1088), .C2(new_n1092), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1106), .B1(new_n1105), .B2(new_n1100), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1096), .B(new_n1142), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT118), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n1096), .A4(new_n1142), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1130), .B1(new_n1144), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(new_n1132), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1108), .B2(new_n1142), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1147), .A2(KEYINPUT118), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n894), .A2(G330), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n273), .A2(new_n857), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n311), .B(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n919), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n913), .B2(new_n918), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1160), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1167), .B2(new_n1165), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1158), .A2(new_n1159), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1132), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1170), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n683), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n827), .B1(new_n202), .B2(new_n796), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n768), .A2(new_n807), .B1(new_n1113), .B2(new_n731), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n752), .B2(G128), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G132), .A2(new_n741), .B1(new_n743), .B2(G137), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(KEYINPUT120), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1179), .B1(new_n1120), .B2(new_n747), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n802), .C2(G159), .ZN(new_n1186));
  INV_X1    g0986(.A(G124), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1187), .B2(new_n758), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT121), .Z(new_n1189));
  NAND3_X1  g0989(.A1(new_n1184), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n802), .A2(G58), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n778), .A2(G283), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n934), .A2(new_n1022), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n742), .B2(new_n504), .C1(new_n356), .C2(new_n744), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n396), .A2(G41), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n747), .B2(new_n219), .C1(new_n363), .C2(new_n751), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1195), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1201));
  AND4_X1   g1001(.A1(new_n1190), .A2(new_n1198), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1177), .B1(new_n815), .B2(new_n1202), .C1(new_n1166), .C2(new_n726), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n1170), .B2(new_n995), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1176), .A2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(new_n1155), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1208), .A2(new_n984), .A3(new_n1142), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n994), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n720), .B1(G68), .B2(new_n797), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n288), .B1(new_n778), .B2(G303), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n336), .B2(new_n735), .C1(new_n504), .C2(new_n731), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n776), .A2(new_n751), .B1(new_n747), .B2(new_n769), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1027), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n363), .B2(new_n744), .C1(new_n219), .C2(new_n742), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1191), .B1(new_n1118), .B2(new_n758), .C1(new_n759), .C2(new_n731), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n408), .B(new_n1217), .C1(G50), .C2(new_n756), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n748), .B1(new_n752), .B2(G137), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n807), .A2(new_n744), .B1(new_n742), .B2(new_n1113), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1216), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1211), .B1(new_n1222), .B2(new_n782), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n850), .B2(new_n726), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1210), .A2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1209), .A2(new_n1225), .ZN(G381));
  NAND3_X1  g1026(.A1(new_n1176), .A2(new_n1153), .A3(new_n1205), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n982), .A2(new_n985), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n994), .B1(new_n1230), .B2(KEYINPUT112), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1229), .B1(new_n1231), .B2(new_n986), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1232), .A2(new_n957), .A3(G390), .ZN(new_n1233));
  OR2_X1    g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(G381), .A2(G384), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1228), .A2(new_n1233), .A3(new_n1235), .ZN(G407));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G343), .C2(new_n1227), .ZN(G409));
  NAND2_X1  g1037(.A1(new_n662), .A2(G213), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1170), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1204), .B1(new_n1240), .B2(new_n985), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(G378), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1173), .A2(new_n984), .A3(new_n1170), .ZN(new_n1243));
  OAI211_X1 g1043(.A(KEYINPUT122), .B(new_n1153), .C1(new_n1243), .C2(new_n1204), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n684), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(new_n1153), .A3(new_n1204), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1238), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1208), .B(KEYINPUT60), .Z(new_n1250));
  NOR2_X1   g1050(.A1(new_n1142), .A2(new_n684), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1225), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1252), .A2(G384), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT123), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1254), .A3(G384), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1252), .B2(G384), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1249), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1249), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n1253), .A3(new_n1255), .A4(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1238), .B(new_n1264), .C1(new_n1245), .C2(new_n1247), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1176), .A2(G378), .A3(new_n1205), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1244), .A3(new_n1242), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1238), .A4(new_n1264), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(new_n1266), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1234), .A2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT124), .ZN(new_n1274));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1017), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(G390), .B1(new_n1232), .B2(new_n957), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(KEYINPUT124), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1017), .A2(new_n1275), .ZN(new_n1282));
  OAI211_X1 g1082(.A(KEYINPUT124), .B(new_n1273), .C1(new_n1233), .C2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1271), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1238), .A4(new_n1264), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1279), .A2(new_n1280), .A3(KEYINPUT61), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1248), .B2(new_n1262), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1265), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1289), .B(new_n1290), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1288), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(G378), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1227), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1287), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1281), .A2(new_n1286), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1227), .A3(new_n1296), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1264), .A2(KEYINPUT126), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT127), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1302), .B(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1306), .A2(new_n1300), .A3(new_n1298), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(G402));
endmodule


