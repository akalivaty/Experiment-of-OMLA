//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT0), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(new_n206), .B2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G13), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n225), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n219), .A2(KEYINPUT1), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n222), .B2(new_n228), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n221), .B(new_n230), .C1(new_n233), .C2(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT65), .Z(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XOR2_X1   g0045(.A(G264), .B(G270), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G58), .B(G77), .Z(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(G77), .A2(new_n257), .B1(new_n263), .B2(G223), .ZN(new_n264));
  INV_X1    g0064(.A(G222), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n258), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT68), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(KEYINPUT68), .A3(new_n273), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G226), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n269), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT71), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n214), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n232), .A2(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n296), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT69), .B1(new_n296), .B2(new_n231), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n272), .B2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n225), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G20), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n302), .C1(G50), .C2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n283), .B2(G169), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n286), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT76), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n305), .A2(KEYINPUT77), .A3(new_n308), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT77), .B1(new_n305), .B2(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n282), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G200), .B2(new_n282), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n310), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n310), .A2(new_n313), .A3(new_n319), .A4(new_n316), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n307), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n294), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n299), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n327));
  OR3_X1    g0127(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n301), .A2(G68), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n256), .A2(G226), .A3(new_n258), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n268), .ZN(new_n335));
  INV_X1    g0135(.A(new_n276), .ZN(new_n336));
  OAI21_X1  g0136(.A(G238), .B1(new_n336), .B2(new_n274), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n281), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT79), .A2(KEYINPUT13), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n339), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n280), .B1(new_n277), .B2(G238), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  OAI21_X1  g0143(.A(G179), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n347), .A3(new_n335), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g0151(.A(KEYINPUT14), .B(new_n345), .C1(new_n346), .C2(new_n348), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n330), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n340), .A2(new_n343), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n330), .B1(new_n354), .B2(G190), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n346), .A2(new_n348), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n356), .A2(KEYINPUT78), .A3(G200), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT78), .B1(new_n356), .B2(G200), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n287), .B(KEYINPUT73), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n232), .A2(new_n323), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n365), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n289), .B(new_n368), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT74), .B(new_n367), .C1(new_n369), .C2(new_n361), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n294), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n366), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n299), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n301), .A2(G77), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n376), .B1(G77), .B2(new_n304), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT75), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n280), .B1(new_n277), .B2(G244), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n263), .A2(G238), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n383));
  INV_X1    g0183(.A(G107), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n383), .C1(new_n384), .C2(new_n256), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n268), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n345), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n379), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n377), .B1(new_n374), .B2(new_n299), .ZN(new_n390));
  INV_X1    g0190(.A(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT75), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n387), .A2(G179), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n293), .B1(new_n272), .B2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(new_n304), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n299), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n293), .A2(new_n398), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(G223), .A2(G1698), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT3), .A2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT3), .A2(G33), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n404), .B1(G226), .B2(new_n258), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G87), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n271), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n271), .A2(new_n273), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n281), .B1(new_n410), .B2(new_n215), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n409), .A2(new_n411), .A3(new_n314), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT7), .B1(new_n256), .B2(G20), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT7), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n261), .A2(new_n418), .A3(new_n232), .A4(new_n262), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(G68), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT80), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G58), .A2(G68), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n232), .B1(new_n234), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n287), .ZN(new_n424));
  INV_X1    g0224(.A(G159), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n421), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n422), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n201), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(KEYINPUT80), .C1(new_n425), .C2(new_n424), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n420), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT16), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT16), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n420), .A2(new_n433), .A3(new_n427), .A4(new_n430), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n299), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n403), .B(new_n416), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n432), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n402), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n412), .B2(new_n284), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT81), .A4(G179), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n443), .A2(new_n444), .B1(G169), .B2(new_n412), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT18), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n412), .A2(G169), .ZN(new_n447));
  INV_X1    g0247(.A(new_n410), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n280), .B1(new_n448), .B2(G232), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n407), .A2(new_n408), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n284), .B(new_n449), .C1(new_n450), .C2(new_n271), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n412), .A2(new_n442), .A3(new_n284), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT18), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(new_n440), .C2(new_n402), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n441), .A2(KEYINPUT17), .A3(new_n416), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n439), .A2(new_n446), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n413), .B1(new_n381), .B2(new_n386), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n387), .A2(new_n314), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n379), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n396), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AND4_X1   g0262(.A1(new_n321), .A2(new_n353), .A3(new_n359), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  OAI211_X1 g0264(.A(G244), .B(new_n258), .C1(new_n405), .C2(new_n406), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n256), .A2(G244), .A3(new_n258), .A4(new_n467), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n466), .A2(KEYINPUT82), .B1(G33), .B2(G283), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n268), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n272), .A2(G45), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(G41), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n480), .A2(G274), .A3(new_n271), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n480), .A2(new_n217), .A3(new_n268), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n474), .A2(G190), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n304), .A2(G97), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n272), .A2(G33), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n304), .B(new_n488), .C1(new_n297), .C2(new_n298), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(new_n216), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n424), .A2(new_n323), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  AND2_X1   g0292(.A1(G97), .A2(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n384), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n491), .B1(new_n497), .B2(G20), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n417), .A2(G107), .A3(new_n419), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n490), .B1(new_n500), .B2(new_n299), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n485), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n483), .B1(new_n473), .B2(new_n268), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n413), .B1(new_n503), .B2(new_n482), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n464), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n474), .A2(new_n482), .A3(new_n484), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G200), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(KEYINPUT83), .A3(new_n501), .A4(new_n485), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n500), .A2(new_n299), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  INV_X1    g0311(.A(new_n490), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n436), .B1(new_n498), .B2(new_n499), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT84), .B1(new_n514), .B2(new_n490), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n474), .A2(G179), .A3(new_n482), .A4(new_n484), .ZN(new_n517));
  AOI211_X1 g0317(.A(new_n483), .B(new_n481), .C1(new_n473), .C2(new_n268), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(new_n345), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT86), .A2(G116), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT86), .A2(G116), .ZN(new_n522));
  OAI21_X1  g0322(.A(G33), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G238), .B(new_n258), .C1(new_n405), .C2(new_n406), .ZN(new_n524));
  OAI211_X1 g0324(.A(G244), .B(G1698), .C1(new_n405), .C2(new_n406), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT85), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n263), .B2(G244), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n268), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G45), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(G1), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n211), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n271), .B1(G274), .B2(new_n531), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G200), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n232), .B1(new_n333), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n494), .A2(new_n210), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n232), .B(G68), .C1(new_n405), .C2(new_n406), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n294), .B2(new_n216), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n299), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n398), .A2(new_n371), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n489), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT87), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(G87), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT87), .B1(new_n489), .B2(new_n210), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n533), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n525), .A2(KEYINPUT85), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n256), .A2(new_n527), .A3(G244), .A4(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n523), .A4(new_n524), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n554), .B2(new_n268), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n535), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n529), .A2(new_n284), .A3(new_n533), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n543), .B(new_n544), .C1(new_n371), .C2(new_n489), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(G169), .C2(new_n555), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n509), .A2(new_n520), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n478), .A2(new_n479), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n268), .B1(new_n531), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n481), .B1(G264), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G294), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n266), .A2(new_n211), .B1(new_n260), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n263), .A2(G257), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(KEYINPUT93), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n314), .B(new_n565), .C1(new_n573), .C2(new_n271), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n564), .A2(G264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n482), .ZN(new_n576));
  INV_X1    g0376(.A(new_n567), .ZN(new_n577));
  INV_X1    g0377(.A(new_n572), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n568), .A2(KEYINPUT93), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n268), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n574), .B1(new_n581), .B2(G200), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n398), .A2(new_n384), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n583), .B(KEYINPUT25), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n489), .A2(new_n384), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT86), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT86), .A2(G116), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n260), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n232), .B2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n384), .A2(KEYINPUT23), .A3(G20), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n591), .A2(new_n232), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT22), .ZN(new_n596));
  AOI21_X1  g0396(.A(G20), .B1(new_n261), .B2(new_n262), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(G87), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n232), .B(G87), .C1(new_n405), .C2(new_n406), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n595), .B(KEYINPUT91), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n256), .A2(new_n596), .A3(new_n232), .A4(G87), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT91), .B1(new_n605), .B2(new_n595), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n595), .B1(new_n598), .B2(new_n600), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT91), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT24), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n299), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n607), .A2(new_n612), .A3(KEYINPUT92), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT92), .ZN(new_n614));
  AOI211_X1 g0414(.A(KEYINPUT91), .B(KEYINPUT24), .C1(new_n605), .C2(new_n595), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n436), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(new_n609), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(KEYINPUT24), .A3(new_n601), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n582), .B(new_n586), .C1(new_n613), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT94), .ZN(new_n621));
  INV_X1    g0421(.A(new_n586), .ZN(new_n622));
  OAI21_X1  g0422(.A(KEYINPUT92), .B1(new_n607), .B2(new_n612), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n618), .A2(new_n614), .A3(new_n299), .A4(new_n611), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT94), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n582), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n562), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n284), .B(new_n565), .C1(new_n573), .C2(new_n271), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n581), .B2(G169), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n586), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n268), .A2(new_n279), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n564), .A2(G270), .B1(new_n633), .B2(new_n480), .ZN(new_n634));
  OAI211_X1 g0434(.A(G264), .B(G1698), .C1(new_n405), .C2(new_n406), .ZN(new_n635));
  OAI211_X1 g0435(.A(G257), .B(new_n258), .C1(new_n405), .C2(new_n406), .ZN(new_n636));
  INV_X1    g0436(.A(G303), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n256), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n268), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n345), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n521), .A2(new_n522), .A3(new_n232), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n296), .A2(new_n231), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT88), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n589), .A2(G20), .A3(new_n590), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT88), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n296), .A2(new_n231), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT20), .ZN(new_n649));
  NAND2_X1  g0449(.A1(G33), .A2(G283), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(new_n232), .C1(G33), .C2(new_n216), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(KEYINPUT89), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n303), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n546), .B2(G116), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n651), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n643), .B2(new_n647), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n649), .A2(KEYINPUT89), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n640), .B1(new_n656), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT21), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT21), .B(new_n640), .C1(new_n656), .C2(new_n662), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n651), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n659), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n660), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(new_n652), .A3(new_n655), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n634), .A2(new_n639), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n284), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n652), .A2(new_n655), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n634), .A2(new_n639), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G190), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n673), .A2(G200), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(new_n678), .A3(new_n671), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n665), .A2(new_n666), .A3(new_n675), .A4(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT90), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n666), .A2(new_n675), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(KEYINPUT90), .A3(new_n665), .A4(new_n680), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n632), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n463), .A2(new_n628), .A3(new_n686), .ZN(G372));
  INV_X1    g0487(.A(KEYINPUT26), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n506), .A2(G169), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n501), .B1(new_n689), .B2(new_n517), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n561), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n557), .A2(new_n516), .A3(new_n519), .A4(new_n560), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n691), .A2(new_n560), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n665), .A2(new_n666), .A3(new_n675), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT95), .B1(new_n632), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n666), .A2(new_n675), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT21), .B1(new_n672), .B2(new_n640), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT95), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n699), .B(new_n700), .C1(new_n625), .C2(new_n630), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n509), .A2(new_n520), .A3(new_n561), .ZN(new_n703));
  AND4_X1   g0503(.A1(new_n626), .A2(new_n631), .A3(new_n586), .A4(new_n582), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n626), .B1(new_n625), .B2(new_n582), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n694), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n463), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT96), .Z(new_n709));
  INV_X1    g0509(.A(new_n353), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n359), .B2(new_n396), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n439), .A2(new_n457), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n446), .B(new_n456), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n318), .A2(new_n320), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n307), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(G369));
  NAND2_X1  g0516(.A1(new_n683), .A2(new_n685), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n653), .A2(KEYINPUT27), .A3(G20), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT27), .B1(new_n653), .B2(G20), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G343), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n672), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n717), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n699), .B2(new_n724), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n632), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n704), .A2(new_n705), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n625), .A2(new_n722), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n632), .A2(new_n722), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n730), .B1(new_n621), .B2(new_n627), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n728), .A3(new_n695), .A4(new_n722), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n732), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(G399));
  INV_X1    g0540(.A(new_n227), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G41), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n538), .A2(G116), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n742), .A2(new_n272), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n236), .B2(new_n742), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  NAND2_X1  g0547(.A1(new_n621), .A2(new_n627), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n748), .A2(new_n696), .A3(new_n703), .A4(new_n701), .ZN(new_n749));
  AOI211_X1 g0549(.A(KEYINPUT29), .B(new_n723), .C1(new_n749), .C2(new_n694), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n699), .B1(new_n625), .B2(new_n630), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n752), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n692), .A2(new_n688), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT97), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT97), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n692), .A2(new_n756), .A3(new_n688), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n690), .A2(KEYINPUT26), .A3(new_n560), .A4(new_n557), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n753), .A2(new_n560), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n751), .B1(new_n760), .B2(new_n722), .ZN(new_n761));
  INV_X1    g0561(.A(G330), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n628), .A2(new_n686), .A3(new_n722), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n581), .A2(new_n503), .A3(new_n555), .A4(new_n674), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT30), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n565), .B1(new_n573), .B2(new_n271), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n677), .A2(G179), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n767), .A2(new_n768), .A3(new_n506), .A4(new_n534), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(new_n764), .B2(new_n765), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n723), .B1(new_n766), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT31), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT31), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n773), .B(new_n723), .C1(new_n766), .C2(new_n770), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n762), .B1(new_n763), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n750), .A2(new_n761), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n747), .B1(new_n777), .B2(G1), .ZN(G364));
  INV_X1    g0578(.A(new_n727), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n225), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n272), .B1(new_n780), .B2(G45), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n742), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G330), .B2(new_n726), .ZN(new_n785));
  INV_X1    g0585(.A(new_n783), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n232), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n413), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n384), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n284), .A2(new_n413), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n787), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n256), .B1(new_n792), .B2(new_n208), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n232), .A2(new_n314), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n284), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n790), .B(new_n793), .C1(G58), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n787), .A2(new_n795), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n323), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n794), .A2(new_n788), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n210), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n791), .A2(new_n794), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n800), .B(new_n802), .C1(G50), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n787), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(KEYINPUT32), .B1(new_n807), .B2(new_n425), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n807), .A2(KEYINPUT32), .A3(new_n425), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n232), .B1(new_n806), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(G97), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n798), .A2(new_n805), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n792), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n814), .A2(new_n815), .B1(new_n797), .B2(G322), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT100), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n257), .B1(new_n799), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G294), .B2(new_n811), .ZN(new_n820));
  INV_X1    g0620(.A(new_n801), .ZN(new_n821));
  INV_X1    g0621(.A(new_n789), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n821), .B1(new_n822), .B2(G283), .ZN(new_n823));
  INV_X1    g0623(.A(new_n807), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n804), .A2(G326), .B1(new_n824), .B2(G329), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n813), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n345), .A2(KEYINPUT99), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n232), .B1(KEYINPUT99), .B2(new_n345), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n231), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n786), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n741), .A2(new_n256), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n530), .B2(new_n236), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n530), .B2(new_n254), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n741), .A2(new_n257), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G355), .B1(new_n588), .B2(new_n741), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(KEYINPUT98), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(KEYINPUT98), .ZN(new_n841));
  NOR2_X1   g0641(.A1(G13), .A2(G33), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(G20), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n844), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n832), .B1(new_n840), .B2(new_n846), .C1(new_n726), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n785), .A2(new_n848), .ZN(G396));
  NAND2_X1  g0649(.A1(new_n707), .A2(new_n722), .ZN(new_n850));
  INV_X1    g0650(.A(new_n461), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n390), .A2(new_n722), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n395), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n392), .A2(new_n389), .A3(new_n394), .A4(new_n852), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n850), .B(new_n856), .Z(new_n857));
  INV_X1    g0657(.A(new_n776), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n783), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n789), .A2(new_n210), .B1(new_n807), .B2(new_n818), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT101), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n589), .A2(new_n590), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n864), .A2(new_n799), .B1(new_n803), .B2(new_n637), .ZN(new_n865));
  INV_X1    g0665(.A(G283), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n384), .A2(new_n801), .B1(new_n792), .B2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n257), .B1(new_n810), .B2(new_n216), .C1(new_n566), .C2(new_n796), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n862), .A2(new_n865), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT102), .ZN(new_n870));
  INV_X1    g0670(.A(G150), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n792), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G143), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n796), .A2(new_n873), .B1(new_n799), .B2(new_n425), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n872), .B(new_n874), .C1(G137), .C2(new_n804), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(KEYINPUT34), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(KEYINPUT34), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n256), .B1(new_n801), .B2(new_n202), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n789), .A2(new_n208), .B1(new_n807), .B2(new_n879), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n878), .B(new_n880), .C1(G58), .C2(new_n811), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n870), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n831), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n831), .A2(new_n842), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n786), .B1(new_n323), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n884), .B(new_n886), .C1(new_n856), .C2(new_n843), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n860), .A2(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n780), .A2(new_n272), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n763), .A2(new_n775), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n463), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT108), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n330), .A2(new_n723), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n359), .A2(new_n353), .A3(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n330), .B(new_n723), .C1(new_n351), .C2(new_n352), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n856), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n763), .B2(new_n775), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n721), .B1(new_n440), .B2(new_n402), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n458), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n454), .B1(new_n440), .B2(new_n402), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n437), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT106), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n903), .A2(new_n437), .A3(new_n907), .A4(new_n900), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n908), .A2(new_n906), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n905), .A2(new_n908), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n902), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n893), .B1(new_n899), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n902), .A2(new_n914), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT40), .B1(new_n920), .B2(new_n915), .ZN(new_n921));
  INV_X1    g0721(.A(new_n898), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n921), .A2(new_n890), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n892), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n892), .A2(new_n924), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(G330), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT109), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n463), .B1(new_n750), .B2(new_n761), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n715), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT107), .Z(new_n932));
  NAND3_X1  g0732(.A1(new_n707), .A2(new_n722), .A3(new_n856), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n395), .A2(new_n723), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT104), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n902), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n902), .B2(new_n914), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n936), .B(new_n897), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n710), .A2(new_n722), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n920), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n937), .B1(new_n911), .B2(new_n912), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(KEYINPUT39), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n446), .A2(new_n456), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n720), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n932), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n889), .B1(new_n929), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n929), .B2(new_n948), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n951), .A2(new_n952), .A3(G116), .A4(new_n233), .ZN(new_n953));
  XOR2_X1   g0753(.A(KEYINPUT103), .B(KEYINPUT36), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n236), .A2(G77), .A3(new_n422), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(G50), .B2(new_n208), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(G1), .A3(new_n225), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n950), .A2(new_n955), .A3(new_n958), .ZN(G367));
  OAI221_X1 g0759(.A(new_n845), .B1(new_n227), .B2(new_n371), .C1(new_n247), .C2(new_n834), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n786), .B1(new_n960), .B2(KEYINPUT114), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT114), .B2(new_n960), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n803), .A2(new_n873), .B1(new_n801), .B2(new_n214), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n257), .B(new_n963), .C1(G150), .C2(new_n797), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n789), .A2(new_n323), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G137), .B2(new_n824), .ZN(new_n966));
  INV_X1    g0766(.A(new_n799), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G159), .A2(new_n814), .B1(new_n967), .B2(G50), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n811), .A2(G68), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n216), .A2(new_n789), .B1(new_n799), .B2(new_n866), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n256), .B(new_n971), .C1(G317), .C2(new_n824), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT115), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT46), .B1(new_n821), .B2(new_n863), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G107), .B2(new_n811), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n803), .A2(new_n818), .B1(new_n796), .B2(new_n637), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(G294), .B2(new_n814), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n972), .A2(new_n974), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n962), .B1(new_n831), .B2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n550), .A2(new_n722), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n561), .A2(new_n983), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n560), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n982), .B1(new_n847), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n781), .B(KEYINPUT113), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n501), .A2(new_n722), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n509), .A2(new_n520), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n690), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n722), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT110), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n509), .A2(new_n520), .A3(new_n990), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n992), .C2(new_n722), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n738), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT112), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n738), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1000), .A2(new_n1002), .A3(KEYINPUT44), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n994), .A2(new_n997), .ZN(new_n1005));
  AOI211_X1 g0805(.A(KEYINPUT112), .B(new_n1005), .C1(new_n737), .C2(new_n732), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1001), .B1(new_n738), .B2(new_n998), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n737), .A2(new_n732), .A3(new_n1005), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n734), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n777), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n699), .A2(new_n723), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n733), .B(new_n1015), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n779), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n733), .B1(new_n699), .B2(new_n723), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n727), .A3(new_n737), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1014), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1003), .A2(new_n1008), .A3(new_n735), .A4(new_n1011), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1013), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n777), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n742), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n989), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n998), .A2(new_n737), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT42), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n520), .B1(new_n998), .B2(new_n728), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n520), .C1(new_n998), .C2(new_n728), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n722), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n986), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT43), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1028), .A2(new_n1033), .A3(new_n1036), .A4(new_n1035), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n735), .A2(new_n998), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1041), .B(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n987), .B1(new_n1026), .B2(new_n1044), .ZN(G387));
  INV_X1    g0845(.A(new_n1020), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1017), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n742), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n293), .A2(new_n792), .B1(new_n208), .B2(new_n799), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT116), .Z(new_n1050));
  NOR2_X1   g0850(.A1(new_n801), .A2(new_n323), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G50), .B2(new_n797), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n804), .A2(G159), .B1(new_n824), .B2(G150), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n810), .A2(new_n371), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n257), .B(new_n1054), .C1(G97), .C2(new_n822), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n256), .B1(new_n824), .B2(G326), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n801), .A2(new_n566), .B1(new_n810), .B2(new_n866), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n792), .A2(new_n818), .ZN(new_n1059));
  INV_X1    g0859(.A(G317), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n796), .A2(new_n1060), .B1(new_n799), .B2(new_n637), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1059), .B(new_n1061), .C1(G322), .C2(new_n804), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1058), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1057), .B1(new_n864), .B2(new_n789), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1056), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n831), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n837), .A2(new_n744), .B1(new_n384), .B2(new_n741), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n369), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n202), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n530), .B1(new_n208), .B2(new_n323), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1073), .A2(new_n744), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n243), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n833), .B1(new_n1076), .B2(new_n530), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n786), .B1(new_n1078), .B2(new_n845), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1069), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n733), .B2(new_n844), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n1082), .B2(new_n989), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1048), .A2(new_n1083), .ZN(G393));
  NAND2_X1  g0884(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1046), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n742), .A3(new_n1022), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT117), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1013), .A2(new_n1021), .A3(new_n989), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n251), .A2(new_n833), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n845), .B1(new_n216), .B2(new_n227), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n783), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n810), .A2(new_n323), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n257), .B(new_n1093), .C1(G87), .C2(new_n822), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n202), .A2(new_n792), .B1(new_n801), .B2(new_n208), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G143), .B2(new_n824), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n369), .C2(new_n799), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n803), .A2(new_n871), .B1(new_n796), .B2(new_n425), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT51), .Z(new_n1099));
  AOI211_X1 g0899(.A(new_n256), .B(new_n790), .C1(new_n863), .C2(new_n811), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G303), .A2(new_n814), .B1(new_n967), .B2(G294), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G283), .A2(new_n821), .B1(new_n824), .B2(G322), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n803), .A2(new_n1060), .B1(new_n796), .B2(new_n818), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT52), .Z(new_n1105));
  OAI22_X1  g0905(.A1(new_n1097), .A2(new_n1099), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1092), .B1(new_n1106), .B2(new_n831), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1005), .B2(new_n847), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n1087), .A2(new_n1088), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1088), .B1(new_n1087), .B2(new_n1110), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(G390));
  AOI21_X1  g0914(.A(new_n786), .B1(new_n293), .B2(new_n885), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G50), .A2(new_n822), .B1(new_n824), .B2(G125), .ZN(new_n1116));
  INV_X1    g0916(.A(G137), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n792), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT53), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n801), .B2(new_n871), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n821), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n256), .B1(new_n799), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n803), .A2(new_n1125), .B1(new_n796), .B2(new_n879), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1124), .B(new_n1126), .C1(G159), .C2(new_n811), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n803), .A2(new_n866), .B1(new_n796), .B2(new_n588), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n792), .A2(new_n384), .B1(new_n807), .B2(new_n566), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n208), .A2(new_n789), .B1(new_n799), .B2(new_n216), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1131), .A2(new_n802), .A3(new_n1093), .A4(new_n256), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1122), .A2(new_n1127), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n831), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1115), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n942), .B1(new_n943), .B2(KEYINPUT39), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n842), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n897), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n933), .B2(new_n935), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1139), .B2(new_n941), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n890), .A2(G330), .A3(new_n856), .A4(new_n897), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n560), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n757), .A2(new_n758), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n755), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n723), .B1(new_n1144), .B2(new_n753), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n934), .B1(new_n1145), .B2(new_n856), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n897), .B(KEYINPUT118), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n916), .B(new_n940), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1140), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1141), .B1(new_n1140), .B2(new_n1148), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1137), .B1(new_n1151), .B2(new_n989), .ZN(new_n1152));
  AND4_X1   g0952(.A1(G330), .A2(new_n890), .A3(new_n856), .A4(new_n897), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n897), .B1(new_n776), .B2(new_n856), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n936), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n890), .A2(G330), .A3(new_n856), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1147), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n1141), .A3(new_n1146), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n463), .A2(new_n776), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n930), .A2(new_n715), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(KEYINPUT119), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1140), .A2(new_n1148), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1153), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n930), .A2(new_n715), .A3(new_n1160), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1140), .A2(new_n1141), .A3(new_n1148), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1163), .A2(new_n742), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT119), .B1(new_n1171), .B2(new_n1162), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1152), .B1(new_n1170), .B2(new_n1172), .ZN(G378));
  NAND2_X1  g0973(.A1(new_n305), .A2(new_n721), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n321), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n321), .A2(new_n1174), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n321), .A2(new_n1174), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1174), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1181), .B(new_n307), .C1(new_n318), .C2(new_n320), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(G330), .C1(new_n917), .C2(new_n923), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n922), .A2(new_n890), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT40), .B1(new_n1187), .B2(new_n943), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n899), .A2(new_n921), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1184), .B1(new_n1190), .B2(G330), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n947), .B1(new_n1186), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1184), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n924), .B2(new_n762), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n947), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n1185), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n786), .B1(new_n202), .B2(new_n885), .ZN(new_n1198));
  INV_X1    g0998(.A(G125), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n803), .A2(new_n1199), .B1(new_n792), .B2(new_n879), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n967), .A2(G137), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n1125), .B2(new_n796), .C1(new_n801), .C2(new_n1123), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G150), .C2(new_n811), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT59), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n822), .A2(G159), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n824), .C2(G124), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1051), .A2(G41), .A3(new_n256), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n822), .A2(G58), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n824), .A2(G283), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n969), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n803), .A2(new_n588), .B1(new_n799), .B2(new_n371), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n216), .A2(new_n792), .B1(new_n796), .B2(new_n384), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n202), .B1(new_n405), .B2(G41), .ZN(new_n1219));
  AND4_X1   g1019(.A1(new_n1209), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1198), .B1(new_n1134), .B2(new_n1220), .C1(new_n1184), .C2(new_n843), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT120), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(KEYINPUT120), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1197), .A2(new_n989), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1169), .A2(new_n1161), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n742), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1197), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1224), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT121), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(KEYINPUT121), .B(new_n1224), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G375));
  AOI21_X1  g1034(.A(new_n786), .B1(new_n208), .B2(new_n885), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n804), .A2(G294), .B1(new_n967), .B2(G107), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n866), .B2(new_n796), .C1(new_n864), .C2(new_n792), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1237), .A2(new_n256), .A3(new_n965), .A4(new_n1054), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n801), .A2(new_n216), .B1(new_n807), .B2(new_n637), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT122), .Z(new_n1240));
  OAI22_X1  g1040(.A1(new_n1117), .A2(new_n796), .B1(new_n801), .B2(new_n425), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n799), .A2(new_n871), .B1(new_n807), .B2(new_n1125), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n803), .A2(new_n879), .B1(new_n792), .B2(new_n1123), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1211), .A2(new_n256), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(G50), .C2(new_n811), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1238), .A2(new_n1240), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1235), .B1(new_n1247), .B2(new_n1134), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1147), .B2(new_n842), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1159), .B2(new_n989), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1162), .A2(new_n1025), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1251), .B2(new_n1252), .ZN(G381));
  NOR3_X1   g1053(.A1(G387), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT123), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT123), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1254), .A2(new_n1258), .A3(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G375), .A2(KEYINPUT125), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1233), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G378), .A2(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT124), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n1152), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1266));
  AND2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1260), .A2(new_n1261), .A3(new_n1263), .A4(new_n1267), .ZN(G407));
  NAND3_X1  g1068(.A1(new_n1261), .A2(new_n1263), .A3(new_n1267), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G343), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(G396), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1022), .A2(new_n742), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1020), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(KEYINPUT117), .B1(new_n1275), .B2(new_n1109), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1087), .A2(new_n1088), .A3(new_n1110), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1041), .B(new_n1042), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1024), .B1(new_n1022), .B2(new_n777), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n989), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1276), .A2(new_n1277), .B1(new_n1280), .B2(new_n987), .ZN(new_n1281));
  OAI211_X1 g1081(.A(KEYINPUT127), .B(new_n1272), .C1(new_n1254), .C2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1272), .A2(KEYINPUT127), .ZN(new_n1283));
  OAI21_X1  g1083(.A(G387), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1276), .A2(new_n1280), .A3(new_n987), .A4(new_n1277), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1272), .A2(KEYINPUT127), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1225), .A2(new_n1197), .A3(new_n1025), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1224), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1264), .A2(new_n1266), .A3(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G378), .B(new_n1224), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(G343), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G213), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G2897), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1166), .A2(new_n1155), .A3(KEYINPUT60), .A4(new_n1158), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n742), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1156), .A2(new_n1138), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1141), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1146), .A2(new_n1141), .ZN(new_n1304));
  AOI22_X1  g1104(.A1(new_n936), .A2(new_n1303), .B1(new_n1304), .B2(new_n1157), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT60), .B1(new_n1305), .B2(new_n1166), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1166), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1301), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1250), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1299), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1252), .B1(KEYINPUT60), .B2(new_n1162), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G384), .B(new_n1250), .C1(new_n1311), .C2(new_n1301), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1298), .B1(new_n1313), .B2(KEYINPUT126), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1298), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1314), .A2(new_n1318), .B1(KEYINPUT126), .B2(new_n1313), .ZN(new_n1319));
  AOI21_X1  g1119(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1295), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1293), .A2(new_n1295), .A3(new_n1313), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1288), .A2(new_n1320), .A3(new_n1323), .A4(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1322), .A2(new_n1328), .A3(new_n1313), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1313), .A2(KEYINPUT126), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1317), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1332));
  AOI211_X1 g1132(.A(KEYINPUT126), .B(new_n1298), .C1(new_n1310), .C2(new_n1312), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1330), .B1(new_n1322), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1328), .B1(new_n1322), .B2(new_n1313), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1329), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1327), .B1(new_n1337), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1138(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1231), .A2(new_n1267), .A3(new_n1232), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(new_n1315), .A3(new_n1292), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1315), .B1(new_n1340), .B2(new_n1292), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1339), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1343), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1345), .A2(new_n1288), .A3(new_n1341), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(G402));
endmodule


