//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G143), .B(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G128), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(G143), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n193), .B(new_n194), .C1(new_n198), .C2(new_n191), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(KEYINPUT0), .A3(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n195), .A2(G143), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n201), .B(new_n202), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n199), .B1(new_n207), .B2(new_n194), .ZN(new_n208));
  INV_X1    g022(.A(G953), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G224), .ZN(new_n210));
  XOR2_X1   g024(.A(new_n210), .B(KEYINPUT81), .Z(new_n211));
  XNOR2_X1  g025(.A(new_n208), .B(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT66), .B1(new_n213), .B2(G116), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(G116), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(KEYINPUT66), .A3(G116), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT2), .A2(G113), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT2), .A2(G113), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n217), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n216), .A2(new_n223), .A3(new_n217), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(G107), .ZN(new_n229));
  INV_X1    g043(.A(G107), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(G104), .C1(KEYINPUT74), .C2(KEYINPUT3), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n228), .A2(G107), .B1(KEYINPUT74), .B2(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n228), .B2(G107), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(G107), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n230), .A2(KEYINPUT75), .A3(G104), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G119), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(G119), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT5), .B(new_n217), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G113), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n246), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT79), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n253), .A3(new_n250), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n225), .A2(new_n242), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n232), .A2(new_n234), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n216), .A2(new_n217), .ZN(new_n262));
  INV_X1    g076(.A(new_n220), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n222), .A2(new_n224), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n255), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(G110), .B(G122), .Z(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT6), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n265), .A2(new_n266), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n265), .A2(KEYINPUT6), .A3(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n212), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n266), .B(new_n276), .Z(new_n277));
  AOI22_X1  g091(.A1(new_n222), .A2(new_n224), .B1(new_n251), .B2(KEYINPUT79), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n242), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n225), .A2(new_n242), .A3(new_n251), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT83), .B(new_n277), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n262), .A2(new_n263), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n225), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n260), .A3(new_n258), .ZN(new_n285));
  INV_X1    g099(.A(new_n266), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n255), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n208), .B(new_n288), .Z(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n225), .A2(new_n254), .A3(new_n252), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n235), .A2(new_n241), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n280), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT83), .B1(new_n294), .B2(new_n277), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n275), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n190), .B1(new_n274), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n212), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n267), .B1(new_n285), .B2(new_n255), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n287), .B1(new_n299), .B2(KEYINPUT6), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n300), .B2(new_n272), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n279), .A2(new_n281), .ZN(new_n303));
  INV_X1    g117(.A(new_n277), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n287), .A3(new_n282), .A4(new_n289), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n301), .A2(new_n306), .A3(new_n275), .A4(new_n189), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n188), .B1(new_n297), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT9), .B(G234), .Z(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n275), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT12), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n197), .B1(new_n196), .B2(KEYINPUT76), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n191), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n192), .A2(G128), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n204), .A2(new_n205), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n235), .B(new_n241), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n191), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n196), .B2(new_n197), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n292), .A2(new_n323), .A3(new_n193), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT11), .ZN(new_n326));
  INV_X1    g140(.A(G134), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G137), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT11), .A3(G134), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n328), .A2(new_n330), .A3(new_n334), .A4(new_n331), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(KEYINPUT64), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n337), .A3(G131), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n313), .B1(new_n325), .B2(new_n340), .ZN(new_n341));
  AOI211_X1 g155(.A(KEYINPUT12), .B(new_n339), .C1(new_n321), .C2(new_n324), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n209), .A2(G227), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT72), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G140), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n346), .B(new_n347), .Z(new_n348));
  NAND3_X1  g162(.A1(new_n258), .A2(new_n207), .A3(new_n260), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n203), .C2(G146), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n317), .A2(G128), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n320), .B1(new_n352), .B2(new_n322), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n353), .B2(new_n292), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n193), .B1(new_n198), .B2(new_n191), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n242), .A2(KEYINPUT10), .A3(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n349), .A2(new_n339), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n343), .A2(new_n344), .A3(new_n348), .A4(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n353), .A2(new_n292), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n355), .B1(new_n235), .B2(new_n241), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n340), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT12), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n325), .A2(new_n313), .A3(new_n340), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n348), .A3(new_n357), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n340), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n357), .ZN(new_n368));
  INV_X1    g182(.A(new_n348), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n275), .ZN(new_n373));
  NAND2_X1  g187(.A1(G469), .A2(G902), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n362), .A2(new_n357), .A3(new_n363), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n348), .B(KEYINPUT73), .Z(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n348), .A3(new_n357), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(G469), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n308), .A2(new_n312), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n336), .A2(new_n207), .A3(new_n338), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT65), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n336), .A2(new_n207), .A3(new_n384), .A4(new_n338), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n327), .A2(G137), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n329), .A2(G134), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n355), .A2(new_n335), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n335), .A2(new_n388), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT68), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(KEYINPUT68), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n355), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(new_n284), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n264), .A3(new_n382), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n209), .A3(G210), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n233), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n402), .B(new_n403), .Z(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT31), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT28), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n390), .A2(new_n284), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n399), .A2(new_n407), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n404), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT31), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n398), .A2(new_n414), .A3(new_n399), .A4(new_n404), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n406), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(G472), .A2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT32), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n396), .A2(new_n382), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n284), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n408), .A2(new_n410), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n404), .A2(KEYINPUT29), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n411), .B2(new_n412), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n404), .B1(new_n398), .B2(new_n399), .ZN(new_n427));
  OAI221_X1 g241(.A(new_n275), .B1(new_n423), .B2(new_n424), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G472), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n416), .A2(KEYINPUT32), .A3(new_n417), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G116), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n230), .B1(new_n434), .B2(KEYINPUT14), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n244), .A2(G122), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n433), .A2(G116), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n244), .A2(G122), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n434), .B(new_n439), .C1(KEYINPUT14), .C2(new_n230), .ZN(new_n440));
  XNOR2_X1  g254(.A(G128), .B(G143), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n327), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n441), .A2(new_n327), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n438), .B(new_n440), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n434), .A2(new_n439), .A3(new_n230), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n230), .B1(new_n434), .B2(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n197), .B2(G143), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n203), .A2(KEYINPUT13), .A3(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n197), .A2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT85), .B1(new_n453), .B2(G134), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(KEYINPUT85), .A3(G134), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT86), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(G134), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G107), .B1(new_n436), .B2(new_n437), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n434), .A2(new_n439), .A3(new_n230), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n461), .A2(new_n462), .B1(new_n327), .B2(new_n441), .ZN(new_n463));
  AND4_X1   g277(.A1(KEYINPUT86), .A2(new_n460), .A3(new_n456), .A4(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n445), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n310), .A2(G217), .A3(new_n209), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n463), .A3(new_n456), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n460), .A2(new_n463), .A3(KEYINPUT86), .A4(new_n456), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n466), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n445), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n432), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n472), .B2(new_n445), .ZN(new_n480));
  INV_X1    g294(.A(new_n445), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n481), .B(new_n466), .C1(new_n470), .C2(new_n471), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n275), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT87), .A3(new_n477), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n275), .B(new_n478), .C1(new_n480), .C2(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n467), .A2(new_n474), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n488), .A2(KEYINPUT88), .A3(new_n275), .A4(new_n478), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n479), .A2(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n228), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n400), .A2(new_n209), .A3(G214), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n203), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G131), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(G143), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n334), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n500));
  INV_X1    g314(.A(G140), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(G125), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(G125), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n194), .A2(G140), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(G146), .B(new_n502), .C1(new_n505), .C2(new_n500), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n502), .B1(new_n505), .B2(new_n500), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n195), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n508), .C1(new_n495), .C2(new_n498), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n499), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n496), .B1(new_n511), .B2(new_n334), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n505), .B(G146), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n512), .B(new_n513), .C1(new_n511), .C2(new_n495), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n492), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n492), .B(new_n514), .C1(new_n499), .C2(new_n509), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n275), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G475), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n209), .A2(G952), .ZN(new_n520));
  INV_X1    g334(.A(G234), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(new_n400), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT21), .B(G898), .Z(new_n523));
  OAI211_X1 g337(.A(G902), .B(G953), .C1(new_n521), .C2(new_n400), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT89), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n505), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT84), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n529), .A2(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(KEYINPUT19), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n528), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n195), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT71), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n506), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n495), .A2(new_n497), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(new_n514), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n516), .B1(new_n539), .B2(new_n492), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n541));
  NOR2_X1   g355(.A1(G475), .A2(G902), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n492), .B1(new_n538), .B2(new_n514), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n517), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n527), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n490), .A2(new_n519), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G110), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n213), .A2(G128), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(G119), .B2(new_n197), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n213), .A2(KEYINPUT23), .A3(G128), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n549), .B(new_n550), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  OR2_X1    g368(.A1(KEYINPUT24), .A2(G110), .ZN(new_n555));
  NAND2_X1  g369(.A1(KEYINPUT24), .A2(G110), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n197), .A2(G119), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n554), .A2(new_n560), .B1(new_n195), .B2(new_n528), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n536), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n550), .A2(new_n558), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n555), .A4(new_n556), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT69), .B1(new_n557), .B2(new_n559), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(G110), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n508), .A2(new_n506), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT70), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT70), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n309), .A2(new_n521), .A3(G953), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n562), .B(new_n575), .C1(new_n570), .C2(new_n571), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G217), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(G234), .B2(new_n275), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(new_n275), .A3(new_n578), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n275), .A4(new_n578), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n584), .B1(new_n589), .B2(new_n581), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n381), .A2(new_n431), .A3(new_n548), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n297), .A2(new_n307), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(new_n187), .A3(new_n526), .A4(new_n590), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n380), .A2(new_n312), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n543), .A2(new_n546), .B1(new_n518), .B2(G475), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n474), .B2(KEYINPUT90), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n488), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(G478), .A3(new_n275), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n483), .A2(new_n476), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n416), .A2(new_n275), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(G472), .B1(new_n416), .B2(new_n417), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n595), .A2(new_n597), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT34), .B(G104), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  NAND3_X1  g423(.A1(new_n543), .A2(new_n546), .A3(KEYINPUT91), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n545), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n519), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n490), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n595), .A2(new_n597), .A3(new_n606), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NAND2_X1  g430(.A1(new_n589), .A2(new_n581), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n572), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n582), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n381), .A2(new_n548), .A3(new_n606), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  OAI21_X1  g438(.A(new_n522), .B1(new_n524), .B2(G900), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n613), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n308), .ZN(new_n627));
  OR3_X1    g441(.A1(new_n626), .A2(new_n627), .A3(KEYINPUT92), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT92), .B1(new_n626), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n621), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n416), .A2(KEYINPUT32), .A3(new_n417), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT32), .B1(new_n416), .B2(new_n417), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n631), .B1(new_n634), .B2(new_n429), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n597), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G128), .ZN(G30));
  NOR4_X1   g452(.A1(new_n621), .A2(new_n188), .A3(new_n490), .A4(new_n598), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT94), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n625), .B(KEYINPUT39), .Z(new_n641));
  NOR2_X1   g455(.A1(new_n596), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT40), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n593), .B(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n640), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n404), .B1(new_n422), .B2(new_n399), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n398), .A2(new_n399), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n404), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n647), .B(new_n652), .C1(KEYINPUT40), .C2(new_n643), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G143), .ZN(G45));
  NAND2_X1  g468(.A1(new_n604), .A2(new_n625), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n627), .A3(new_n596), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n635), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G146), .ZN(G48));
  INV_X1    g472(.A(new_n590), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n634), .B2(new_n429), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n371), .A2(new_n275), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G469), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT95), .A3(new_n373), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT95), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n664), .A3(G469), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n311), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n604), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n668), .A2(new_n627), .A3(new_n527), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT41), .B(G113), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G15));
  AND3_X1   g486(.A1(new_n613), .A2(new_n308), .A3(new_n526), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G116), .ZN(G18));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n308), .A3(new_n548), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n431), .A2(new_n621), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n213), .ZN(G21));
  NAND2_X1  g493(.A1(new_n479), .A2(new_n484), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n487), .A2(new_n489), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n543), .A2(new_n546), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n519), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT96), .B1(new_n490), .B2(new_n598), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n308), .A2(new_n686), .A3(new_n687), .A4(new_n526), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n423), .A2(new_n412), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n406), .A2(new_n415), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n417), .ZN(new_n691));
  INV_X1    g505(.A(G472), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n416), .B2(new_n275), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n691), .A2(new_n693), .A3(new_n659), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n688), .A2(new_n666), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  NAND2_X1  g510(.A1(new_n663), .A2(new_n665), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n308), .A3(new_n312), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n655), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n631), .A2(new_n691), .A3(new_n693), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  NAND3_X1  g517(.A1(new_n297), .A2(new_n307), .A3(new_n187), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT97), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n377), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n375), .A2(KEYINPUT97), .A3(new_n376), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n378), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n373), .B(new_n374), .C1(new_n709), .C2(new_n372), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n705), .A2(new_n312), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n660), .A2(new_n700), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n710), .A2(new_n312), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n431), .A2(new_n715), .A3(new_n590), .A4(new_n705), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  INV_X1    g533(.A(new_n626), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n660), .A2(new_n720), .A3(new_n711), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT98), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT98), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n716), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  AND2_X1   g540(.A1(new_n602), .A2(new_n603), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n685), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT43), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT99), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n605), .A2(G472), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n418), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n728), .A2(KEYINPUT43), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT99), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(KEYINPUT43), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n730), .A2(new_n732), .A3(new_n621), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n377), .A2(new_n378), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n372), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n709), .B2(new_n741), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(new_n374), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  INV_X1    g559(.A(new_n373), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n311), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n641), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n705), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n737), .B2(new_n738), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G137), .ZN(G39));
  XNOR2_X1  g567(.A(new_n748), .B(KEYINPUT47), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n431), .A2(new_n655), .A3(new_n590), .A4(new_n704), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT100), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n754), .A2(KEYINPUT100), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n666), .A2(new_n705), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n765), .B(new_n522), .C1(new_n733), .C2(new_n735), .ZN(new_n766));
  INV_X1    g580(.A(new_n522), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT107), .B1(new_n729), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(KEYINPUT112), .B(new_n764), .C1(new_n766), .C2(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n762), .B1(new_n773), .B2(new_n701), .ZN(new_n774));
  INV_X1    g588(.A(new_n701), .ZN(new_n775));
  AOI211_X1 g589(.A(KEYINPUT113), .B(new_n775), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT111), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n694), .B1(new_n766), .B2(new_n768), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n666), .A2(new_n188), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n646), .B1(new_n781), .B2(KEYINPUT109), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(KEYINPUT109), .B2(new_n781), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n780), .B1(KEYINPUT110), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n783), .A2(KEYINPUT110), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n779), .A3(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n652), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n764), .A2(new_n767), .A3(new_n590), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n727), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n685), .A3(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n694), .B(new_n705), .C1(new_n766), .C2(new_n768), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n697), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n798), .A3(new_n312), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n754), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n777), .A2(new_n789), .A3(KEYINPUT51), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n801), .B1(new_n774), .B2(new_n776), .ZN(new_n804));
  INV_X1    g618(.A(new_n788), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n786), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OAI221_X1 g621(.A(new_n520), .B1(new_n668), .B2(new_n791), .C1(new_n780), .C2(new_n698), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n773), .A2(new_n660), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n802), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n695), .A2(new_n607), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n699), .A2(new_n548), .A3(new_n635), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n660), .B(new_n666), .C1(new_n669), .C2(new_n673), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n591), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n490), .A2(new_n685), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n595), .A2(new_n597), .A3(new_n606), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT101), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n622), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n622), .B2(new_n820), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT102), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n714), .A2(new_n717), .B1(new_n722), .B2(new_n724), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n490), .A2(new_n519), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n610), .A2(new_n611), .A3(new_n625), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n704), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n635), .A2(new_n597), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n711), .A2(new_n700), .A3(new_n701), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n819), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n732), .A2(new_n594), .A3(new_n596), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n548), .A2(new_n308), .A3(new_n312), .A4(new_n380), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n732), .A3(new_n631), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT101), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n622), .A2(new_n820), .A3(new_n821), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n695), .A2(new_n591), .A3(new_n607), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n678), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n843), .A3(new_n817), .A4(new_n833), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n718), .A2(new_n725), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT102), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n686), .A2(new_n687), .A3(new_n308), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n631), .A2(new_n625), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n652), .A2(new_n848), .A3(new_n715), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT103), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n850), .B(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n702), .B(new_n657), .C1(new_n636), .C2(new_n630), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n850), .B(KEYINPUT103), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n775), .A2(new_n655), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n856), .A2(new_n699), .B1(new_n635), .B2(new_n656), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(KEYINPUT52), .A3(new_n637), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n834), .A2(new_n846), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT104), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(new_n859), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n834), .A2(new_n846), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n862), .A2(new_n863), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n844), .A2(new_n845), .A3(new_n861), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n865), .B(new_n874), .C1(new_n866), .C2(new_n859), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n860), .A2(KEYINPUT106), .A3(new_n861), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT106), .B1(new_n860), .B2(new_n861), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n814), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n814), .A2(new_n872), .A3(KEYINPUT115), .A4(new_n878), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT116), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n728), .A2(new_n187), .A3(new_n312), .A4(new_n590), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n646), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n796), .A2(KEYINPUT49), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n790), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n209), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT56), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(G902), .ZN(new_n896));
  INV_X1    g710(.A(G210), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n271), .A2(new_n273), .A3(new_n212), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n301), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n893), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n898), .B2(new_n901), .ZN(G51));
  NOR2_X1   g717(.A1(new_n896), .A2(new_n743), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n374), .B(KEYINPUT57), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n860), .A2(new_n861), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT106), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n860), .A2(KEYINPUT106), .A3(new_n861), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n873), .B1(new_n910), .B2(new_n875), .ZN(new_n911));
  INV_X1    g725(.A(new_n878), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n371), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n914), .B2(KEYINPUT117), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n916), .A3(new_n371), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n892), .B1(new_n915), .B2(new_n917), .ZN(G54));
  AND2_X1   g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n895), .A2(G902), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n540), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n892), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n895), .A2(G902), .A3(new_n540), .A4(new_n919), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(KEYINPUT118), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT119), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n928), .B(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(new_n872), .A2(new_n878), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT59), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n601), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n911), .A2(new_n912), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n601), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n893), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT60), .Z(new_n940));
  NAND3_X1  g754(.A1(new_n895), .A2(new_n619), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n895), .A2(new_n940), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(KEYINPUT121), .A3(new_n579), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n579), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n945), .A2(new_n947), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n949), .A2(new_n893), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n944), .B2(new_n943), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n952), .B1(KEYINPUT61), .B2(new_n954), .ZN(G66));
  AOI21_X1  g769(.A(new_n209), .B1(new_n523), .B2(G224), .ZN(new_n956));
  INV_X1    g770(.A(new_n825), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n209), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n271), .B(new_n273), .C1(G898), .C2(new_n209), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(G69));
  OR2_X1    g774(.A1(new_n853), .A2(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n853), .A2(KEYINPUT122), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n653), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n760), .A2(new_n752), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n704), .B1(new_n668), .B2(new_n835), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n660), .A2(new_n642), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT123), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n965), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n392), .A2(new_n397), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n533), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n209), .A3(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(G227), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n209), .B1(new_n979), .B2(G900), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n748), .A2(new_n660), .A3(new_n749), .A4(new_n848), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n961), .A2(new_n962), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n827), .B(KEYINPUT124), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n966), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n209), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n978), .B2(G953), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n980), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n977), .A2(new_n987), .ZN(G72));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n984), .B2(new_n957), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n649), .B(KEYINPUT125), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(new_n412), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n892), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n971), .A2(new_n825), .A3(new_n973), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n990), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n992), .A2(new_n412), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n998), .ZN(new_n1000));
  AOI211_X1 g814(.A(KEYINPUT126), .B(new_n1000), .C1(new_n996), .C2(new_n990), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n994), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n427), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n405), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n990), .B(new_n1004), .C1(new_n870), .C2(new_n871), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1002), .A2(new_n1007), .ZN(G57));
endmodule


