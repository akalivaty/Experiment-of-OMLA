

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  NAND2_X1 U320 ( .A1(G230GAT), .A2(G233GAT), .ZN(n288) );
  NAND2_X1 U321 ( .A1(n375), .A2(n476), .ZN(n376) );
  NOR2_X1 U322 ( .A1(n377), .A2(n376), .ZN(n379) );
  XNOR2_X1 U323 ( .A(n330), .B(n288), .ZN(n331) );
  XNOR2_X1 U324 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n387) );
  XNOR2_X1 U325 ( .A(n332), .B(n331), .ZN(n334) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n520) );
  INV_X1 U327 ( .A(G190GAT), .ZN(n442) );
  NOR2_X1 U328 ( .A1(n522), .A2(n441), .ZN(n556) );
  XOR2_X1 U329 ( .A(n460), .B(KEYINPUT28), .Z(n524) );
  XNOR2_X1 U330 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U331 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G120GAT), .B(G71GAT), .Z(n325) );
  XOR2_X1 U333 ( .A(KEYINPUT85), .B(G190GAT), .Z(n290) );
  XNOR2_X1 U334 ( .A(G15GAT), .B(G99GAT), .ZN(n289) );
  XNOR2_X1 U335 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U336 ( .A(n325), .B(n291), .Z(n293) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(G43GAT), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U339 ( .A(G127GAT), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n416) );
  XOR2_X1 U342 ( .A(G176GAT), .B(n416), .Z(n297) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U346 ( .A(KEYINPUT17), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT19), .B(n302), .ZN(n400) );
  XOR2_X1 U350 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT84), .B(KEYINPUT65), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U353 ( .A(n400), .B(n305), .Z(n306) );
  XOR2_X1 U354 ( .A(n307), .B(n306), .Z(n512) );
  INV_X1 U355 ( .A(n512), .ZN(n522) );
  XOR2_X1 U356 ( .A(KEYINPUT69), .B(KEYINPUT7), .Z(n309) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT8), .B(n310), .Z(n352) );
  XOR2_X1 U360 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n312) );
  XNOR2_X1 U361 ( .A(G113GAT), .B(KEYINPUT67), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n352), .B(n313), .ZN(n324) );
  XOR2_X1 U364 ( .A(G169GAT), .B(G8GAT), .Z(n397) );
  XOR2_X1 U365 ( .A(G197GAT), .B(G141GAT), .Z(n315) );
  XNOR2_X1 U366 ( .A(G36GAT), .B(G50GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(n397), .B(n316), .Z(n318) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n319), .B(KEYINPUT68), .Z(n322) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G15GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n320), .B(G1GAT), .ZN(n369) );
  XNOR2_X1 U374 ( .A(n369), .B(KEYINPUT29), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n492) );
  INV_X1 U377 ( .A(n492), .ZN(n563) );
  XOR2_X1 U378 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n327) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .Z(n370) );
  XNOR2_X1 U380 ( .A(n325), .B(n370), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n332) );
  XOR2_X1 U382 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n329) );
  XNOR2_X1 U383 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G204GAT), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(G64GAT), .ZN(n389) );
  XNOR2_X1 U387 ( .A(n334), .B(n389), .ZN(n340) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(G78GAT), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(G148GAT), .ZN(n431) );
  XOR2_X1 U390 ( .A(KEYINPUT72), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(KEYINPUT73), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U393 ( .A(G85GAT), .B(n338), .Z(n344) );
  XNOR2_X1 U394 ( .A(n431), .B(n344), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n568) );
  XNOR2_X1 U396 ( .A(n568), .B(KEYINPUT41), .ZN(n540) );
  NAND2_X1 U397 ( .A1(n563), .A2(n540), .ZN(n341) );
  XOR2_X1 U398 ( .A(KEYINPUT46), .B(n341), .Z(n377) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n343) );
  XOR2_X1 U400 ( .A(G50GAT), .B(G162GAT), .Z(n426) );
  XOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .Z(n392) );
  XNOR2_X1 U402 ( .A(n426), .B(n392), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U404 ( .A(n345), .B(n344), .Z(n347) );
  XNOR2_X1 U405 ( .A(G218GAT), .B(G106GAT), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U407 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n349) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U410 ( .A(n351), .B(n350), .Z(n354) );
  XNOR2_X1 U411 ( .A(n352), .B(G134GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n545) );
  INV_X1 U413 ( .A(n545), .ZN(n375) );
  XOR2_X1 U414 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n356) );
  XNOR2_X1 U415 ( .A(KEYINPUT80), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n368) );
  XOR2_X1 U417 ( .A(G78GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U418 ( .A(G183GAT), .B(G211GAT), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n366) );
  XOR2_X1 U420 ( .A(KEYINPUT81), .B(KEYINPUT78), .Z(n360) );
  XNOR2_X1 U421 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G71GAT), .Z(n362) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(G127GAT), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U426 ( .A(n364), .B(n363), .Z(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n374) );
  XOR2_X1 U429 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n572) );
  INV_X1 U433 ( .A(n572), .ZN(n476) );
  INV_X1 U434 ( .A(KEYINPUT47), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n386) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(n545), .Z(n578) );
  NOR2_X1 U437 ( .A1(n578), .A2(n476), .ZN(n382) );
  XOR2_X1 U438 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n380) );
  XNOR2_X1 U439 ( .A(KEYINPUT66), .B(n380), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n383) );
  NAND2_X1 U441 ( .A1(n568), .A2(n383), .ZN(n384) );
  NOR2_X1 U442 ( .A1(n384), .A2(n563), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n386), .A2(n385), .ZN(n388) );
  XOR2_X1 U444 ( .A(n389), .B(G92GAT), .Z(n391) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U447 ( .A(n393), .B(n392), .Z(n399) );
  XOR2_X1 U448 ( .A(KEYINPUT21), .B(G218GAT), .Z(n395) );
  XNOR2_X1 U449 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U451 ( .A(G197GAT), .B(n396), .Z(n434) );
  XNOR2_X1 U452 ( .A(n397), .B(n434), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n402) );
  INV_X1 U454 ( .A(n400), .ZN(n401) );
  XOR2_X1 U455 ( .A(n402), .B(n401), .Z(n450) );
  OR2_X1 U456 ( .A1(n520), .A2(n450), .ZN(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT54), .B(n403), .ZN(n558) );
  XOR2_X1 U458 ( .A(KEYINPUT90), .B(G148GAT), .Z(n405) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G120GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U461 ( .A(G162GAT), .B(G85GAT), .Z(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n420) );
  XOR2_X1 U463 ( .A(G57GAT), .B(KEYINPUT4), .Z(n409) );
  XNOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U466 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n411) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U469 ( .A(n413), .B(n412), .Z(n418) );
  XOR2_X1 U470 ( .A(G155GAT), .B(KEYINPUT2), .Z(n415) );
  XNOR2_X1 U471 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n433) );
  XNOR2_X1 U473 ( .A(n416), .B(n433), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n422) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n457) );
  XOR2_X1 U478 ( .A(G204GAT), .B(KEYINPUT86), .Z(n424) );
  XNOR2_X1 U479 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U481 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n438) );
  XOR2_X1 U484 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n430) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U490 ( .A(n438), .B(n437), .Z(n460) );
  NAND2_X1 U491 ( .A1(n457), .A2(n460), .ZN(n439) );
  NOR2_X1 U492 ( .A1(n558), .A2(n439), .ZN(n440) );
  XNOR2_X1 U493 ( .A(KEYINPUT55), .B(n440), .ZN(n441) );
  NAND2_X1 U494 ( .A1(n556), .A2(n545), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT34), .B(KEYINPUT97), .Z(n466) );
  NAND2_X1 U497 ( .A1(n563), .A2(n568), .ZN(n479) );
  NOR2_X1 U498 ( .A1(n545), .A2(n476), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT16), .ZN(n464) );
  NOR2_X1 U500 ( .A1(n460), .A2(n512), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT95), .B(n447), .Z(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT26), .B(n448), .Z(n537) );
  INV_X1 U503 ( .A(n537), .ZN(n560) );
  INV_X1 U504 ( .A(n450), .ZN(n509) );
  XOR2_X1 U505 ( .A(n509), .B(KEYINPUT93), .Z(n449) );
  XNOR2_X1 U506 ( .A(n449), .B(KEYINPUT27), .ZN(n458) );
  NAND2_X1 U507 ( .A1(n560), .A2(n458), .ZN(n455) );
  NOR2_X1 U508 ( .A1(n522), .A2(n450), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT96), .B(n451), .Z(n452) );
  NAND2_X1 U510 ( .A1(n460), .A2(n452), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT25), .B(n453), .Z(n454) );
  NAND2_X1 U512 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n456), .A2(n457), .ZN(n463) );
  INV_X1 U514 ( .A(n457), .ZN(n559) );
  NAND2_X1 U515 ( .A1(n458), .A2(n559), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT94), .ZN(n519) );
  NOR2_X1 U517 ( .A1(n519), .A2(n524), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n522), .A2(n461), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n475) );
  NAND2_X1 U520 ( .A1(n464), .A2(n475), .ZN(n493) );
  NOR2_X1 U521 ( .A1(n479), .A2(n493), .ZN(n472) );
  NAND2_X1 U522 ( .A1(n472), .A2(n559), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  NAND2_X1 U525 ( .A1(n509), .A2(n472), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n468), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n470) );
  NAND2_X1 U528 ( .A1(n472), .A2(n512), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U530 ( .A(G15GAT), .B(n471), .ZN(G1326GAT) );
  XOR2_X1 U531 ( .A(G22GAT), .B(KEYINPUT99), .Z(n474) );
  NAND2_X1 U532 ( .A1(n472), .A2(n524), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1327GAT) );
  XOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT39), .Z(n483) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n477), .A2(n578), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT37), .ZN(n504) );
  NOR2_X1 U538 ( .A1(n504), .A2(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n489) );
  NAND2_X1 U541 ( .A1(n489), .A2(n559), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  NAND2_X1 U543 ( .A1(n489), .A2(n509), .ZN(n484) );
  XNOR2_X1 U544 ( .A(G36GAT), .B(n484), .ZN(G1329GAT) );
  XNOR2_X1 U545 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n486) );
  NAND2_X1 U547 ( .A1(n489), .A2(n512), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1330GAT) );
  XOR2_X1 U550 ( .A(G50GAT), .B(KEYINPUT103), .Z(n491) );
  NAND2_X1 U551 ( .A1(n489), .A2(n524), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1331GAT) );
  XNOR2_X1 U553 ( .A(KEYINPUT104), .B(n540), .ZN(n553) );
  NAND2_X1 U554 ( .A1(n553), .A2(n492), .ZN(n505) );
  NOR2_X1 U555 ( .A1(n505), .A2(n493), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT105), .B(n494), .Z(n500) );
  NAND2_X1 U557 ( .A1(n500), .A2(n559), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(KEYINPUT42), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(n496), .ZN(G1332GAT) );
  NAND2_X1 U560 ( .A1(n509), .A2(n500), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U562 ( .A(G64GAT), .B(n498), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n512), .A2(n500), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n499), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n502) );
  NAND2_X1 U566 ( .A1(n500), .A2(n524), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U568 ( .A(G78GAT), .B(n503), .Z(G1335GAT) );
  XOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT109), .Z(n508) );
  NOR2_X1 U570 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT108), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n559), .A2(n515), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n509), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(KEYINPUT110), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(n511), .ZN(G1337GAT) );
  XOR2_X1 U577 ( .A(G99GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U578 ( .A1(n515), .A2(n512), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n517) );
  NAND2_X1 U581 ( .A1(n524), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n518), .Z(G1339GAT) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n521), .Z(n538) );
  NOR2_X1 U587 ( .A1(n522), .A2(n538), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT115), .B(n523), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n563), .A2(n534), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U593 ( .A1(n534), .A2(n553), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n531) );
  NAND2_X1 U597 ( .A1(n534), .A2(n572), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U601 ( .A1(n534), .A2(n545), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n563), .A2(n546), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  NAND2_X1 U607 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n572), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U612 ( .A(G162GAT), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n556), .A2(n563), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n551) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT120), .B(n552), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n556), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n572), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  AND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT123), .B(n562), .ZN(n577) );
  INV_X1 U628 ( .A(n577), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n573), .A2(n563), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n565) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XNOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n570) );
  NOR2_X1 U635 ( .A1(n577), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(G204GAT), .B(n571), .Z(G1353GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n576) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

