//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(G238), .Z(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT67), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n210), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n212), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n232), .B(new_n235), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n226), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT17), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT78), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT69), .A2(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT69), .A2(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(G68), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n210), .B1(new_n257), .B2(new_n227), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G159), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n254), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(G20), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(KEYINPUT7), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT7), .ZN(new_n269));
  AOI211_X1 g0069(.A(new_n269), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n270));
  OAI21_X1  g0070(.A(G68), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT69), .B(G58), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n201), .B1(new_n272), .B2(G68), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT78), .B(new_n260), .C1(new_n273), .C2(new_n210), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n262), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n264), .A2(new_n266), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(KEYINPUT77), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n269), .B1(new_n280), .B2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT77), .B1(new_n267), .B2(KEYINPUT7), .ZN(new_n283));
  OAI21_X1  g0083(.A(G68), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(KEYINPUT16), .A3(new_n262), .A4(new_n274), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n211), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n230), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n277), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  OAI21_X1  g0089(.A(G58), .B1(new_n289), .B2(KEYINPUT8), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n289), .B2(KEYINPUT8), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT8), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT70), .B1(new_n272), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n255), .A2(new_n256), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT8), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n291), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g0099(.A1(G1), .A2(G13), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n211), .B2(G33), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G1), .B2(new_n210), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n299), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n288), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT68), .B(G41), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  AOI21_X1  g0107(.A(G1), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n309));
  INV_X1    g0109(.A(G274), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G41), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n307), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G41), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n209), .A2(new_n313), .B1(new_n300), .B2(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n308), .A2(new_n311), .B1(G232), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n264), .A2(new_n266), .A3(G226), .A4(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n264), .A2(new_n266), .A3(G223), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G33), .A2(G87), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n309), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(G190), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(KEYINPUT79), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT79), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n253), .B1(new_n305), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n316), .A2(new_n322), .A3(new_n326), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n326), .B1(new_n316), .B2(new_n322), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n334), .B1(G190), .B2(new_n323), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(KEYINPUT17), .A3(new_n304), .A4(new_n288), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n331), .A2(KEYINPUT80), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT18), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n323), .A2(G179), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n328), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n305), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n305), .A2(new_n338), .A3(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT80), .B1(new_n331), .B2(new_n336), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n337), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n308), .A2(new_n311), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G226), .B2(new_n315), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n280), .A2(G223), .A3(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n280), .A2(new_n318), .ZN(new_n352));
  INV_X1    g0152(.A(G222), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n350), .B1(new_n351), .B2(new_n280), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n309), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n340), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G179), .B2(new_n356), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n210), .A2(G33), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n297), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n287), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n298), .A2(G50), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n303), .B2(G50), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(KEYINPUT73), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n365), .A2(KEYINPUT9), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n365), .A2(KEYINPUT9), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n368), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n367), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n302), .A2(new_n216), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT74), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n351), .B2(new_n360), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n381), .A2(new_n287), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(KEYINPUT11), .ZN(new_n383));
  INV_X1    g0183(.A(new_n298), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n216), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n382), .A2(KEYINPUT11), .ZN(new_n387));
  AND4_X1   g0187(.A1(new_n379), .A2(new_n383), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n352), .C2(new_n214), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n309), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n308), .A2(new_n311), .B1(G238), .B2(new_n315), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n388), .B1(new_n369), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n329), .B1(new_n395), .B2(new_n397), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(G169), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G179), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n340), .B1(new_n395), .B2(new_n397), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT76), .A3(new_n402), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT14), .B1(new_n410), .B2(KEYINPUT75), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n398), .A2(KEYINPUT75), .A3(G169), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n409), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n388), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n401), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT8), .B(G58), .ZN(new_n417));
  INV_X1    g0217(.A(new_n259), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n210), .B2(new_n351), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(new_n360), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n287), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n384), .A2(new_n351), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n351), .C2(new_n302), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n348), .B1(G244), .B2(new_n315), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n280), .A2(G232), .A3(new_n318), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n280), .A2(G1698), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n428), .B1(new_n206), .B2(new_n280), .C1(new_n429), .C2(new_n215), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n309), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n425), .A2(new_n426), .B1(new_n432), .B2(new_n369), .ZN(new_n433));
  INV_X1    g0233(.A(new_n432), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n329), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n406), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n340), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n438), .A2(new_n424), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n436), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AND4_X1   g0240(.A1(new_n347), .A2(new_n377), .A3(new_n416), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n259), .A2(G77), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT6), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n446), .A2(new_n205), .A3(G107), .ZN(new_n447));
  XNOR2_X1  g0247(.A(G97), .B(G107), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n445), .B1(new_n210), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n267), .A2(KEYINPUT7), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n206), .B1(new_n451), .B2(new_n281), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n287), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n298), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n209), .A2(G33), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n301), .A2(new_n298), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(G97), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n300), .A2(new_n314), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n209), .B(G45), .C1(new_n463), .C2(G41), .ZN(new_n464));
  OAI211_X1 g0264(.A(G257), .B(new_n461), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n312), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G41), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n464), .B1(new_n469), .B2(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n311), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n280), .A2(G244), .A3(new_n318), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT4), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n318), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n479), .B2(new_n309), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G190), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n460), .B(new_n481), .C1(new_n329), .C2(new_n480), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n280), .A2(new_n210), .A3(G68), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n210), .B1(new_n390), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(G87), .B2(new_n207), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n360), .B2(new_n205), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n488), .A2(new_n287), .B1(new_n384), .B2(new_n420), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n457), .A2(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n280), .A2(G244), .A3(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n280), .A2(G238), .A3(new_n318), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n493), .B(new_n494), .C1(new_n263), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n309), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n209), .A2(new_n310), .A3(G45), .ZN(new_n498));
  INV_X1    g0298(.A(G250), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n307), .B2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n461), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  INV_X1    g0303(.A(new_n501), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n496), .B2(new_n309), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .A3(G190), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT82), .B1(new_n505), .B2(G190), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n492), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(new_n309), .ZN(new_n510));
  INV_X1    g0310(.A(new_n472), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n510), .A2(new_n511), .A3(G179), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n340), .B1(new_n510), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n459), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n489), .B1(new_n420), .B2(new_n456), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n505), .A2(new_n406), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(G169), .C2(new_n505), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n482), .A2(new_n509), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n206), .A2(G20), .ZN(new_n520));
  OAI22_X1  g0320(.A1(KEYINPUT23), .A2(new_n520), .B1(new_n360), .B2(new_n495), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT86), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n520), .B2(KEYINPUT23), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n520), .A2(new_n522), .A3(KEYINPUT23), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n280), .A2(new_n528), .A3(new_n210), .A4(G87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n280), .A2(new_n210), .A3(G87), .ZN(new_n530));
  INV_X1    g0330(.A(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n526), .A2(new_n527), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n524), .A3(new_n529), .A4(new_n525), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n301), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n384), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT25), .B1(new_n384), .B2(new_n206), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n456), .A2(new_n206), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n280), .A2(G257), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n352), .C2(new_n499), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n470), .A2(new_n309), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n309), .A2(new_n544), .B1(new_n545), .B2(G264), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(G190), .A3(new_n471), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n471), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n541), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n340), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n406), .A3(new_n471), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n536), .C2(new_n540), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n502), .B2(new_n369), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n506), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n491), .B1(G200), .B2(new_n502), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n505), .A2(new_n406), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n505), .A2(G169), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n558), .A2(new_n559), .B1(new_n562), .B2(new_n515), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT83), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n514), .A4(new_n482), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n478), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n495), .A2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n287), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n287), .A2(KEYINPUT20), .A3(new_n566), .A4(new_n567), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(KEYINPUT84), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n298), .A2(new_n495), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n457), .B2(new_n495), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT84), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n568), .A2(new_n575), .A3(new_n569), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n280), .A2(G257), .A3(new_n318), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  INV_X1    g0379(.A(G264), .ZN(new_n580));
  OAI221_X1 g0380(.A(new_n578), .B1(new_n579), .B2(new_n280), .C1(new_n429), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n309), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n545), .A2(G270), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n471), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n577), .A2(G169), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(G200), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n369), .C2(new_n584), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n582), .A2(G179), .A3(new_n471), .A4(new_n583), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n577), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n577), .A2(KEYINPUT21), .A3(G169), .A4(new_n584), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n587), .A2(new_n590), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n519), .A2(new_n555), .A3(new_n565), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n442), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0398(.A(new_n344), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n342), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n437), .A2(new_n424), .A3(new_n438), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT89), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n439), .A2(KEYINPUT89), .A3(new_n437), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n401), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n415), .B2(new_n414), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n337), .A2(new_n346), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n600), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n375), .A2(new_n376), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n367), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n512), .A2(new_n513), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT88), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n509), .A2(new_n459), .A3(new_n517), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n512), .A2(new_n513), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(new_n509), .A3(new_n459), .A4(new_n517), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n619), .A2(KEYINPUT26), .B1(new_n515), .B2(new_n562), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n593), .A2(new_n594), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n587), .ZN(new_n622));
  INV_X1    g0422(.A(new_n553), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n563), .A2(new_n550), .A3(new_n514), .A4(new_n482), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n617), .B(new_n620), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n612), .B1(new_n442), .B2(new_n627), .ZN(G369));
  NAND3_X1  g0428(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(G343), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n577), .A2(new_n634), .ZN(new_n635));
  MUX2_X1   g0435(.A(new_n622), .B(new_n595), .S(new_n635), .Z(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(G330), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n553), .A2(new_n634), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n548), .A2(new_n369), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n329), .B1(new_n546), .B2(new_n471), .ZN(new_n641));
  NOR4_X1   g0441(.A1(new_n640), .A2(new_n536), .A3(new_n641), .A4(new_n540), .ZN(new_n642));
  INV_X1    g0442(.A(new_n634), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n541), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n639), .B1(new_n645), .B2(new_n623), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n637), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n634), .B1(new_n621), .B2(new_n587), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n639), .A3(new_n650), .ZN(G399));
  NAND2_X1  g0451(.A1(new_n233), .A2(new_n306), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n228), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n517), .B(KEYINPUT90), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n619), .B2(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n614), .A2(new_n615), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(KEYINPUT26), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT91), .B1(new_n622), .B2(new_n623), .ZN(new_n662));
  INV_X1    g0462(.A(new_n625), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n621), .A2(new_n664), .A3(new_n553), .A4(new_n587), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n657), .B1(new_n667), .B2(new_n643), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n626), .A2(new_n657), .A3(new_n643), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G330), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n554), .B1(new_n518), .B2(KEYINPUT83), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n595), .A3(new_n565), .A4(new_n643), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n546), .A2(new_n505), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n592), .A2(KEYINPUT30), .A3(new_n674), .A4(new_n480), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n546), .A2(new_n510), .A3(new_n511), .A4(new_n505), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n591), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n510), .A2(new_n511), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n505), .A2(G179), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n679), .A2(new_n548), .A3(new_n584), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n634), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT31), .B1(new_n682), .B2(new_n634), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n671), .B1(new_n673), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n670), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n656), .B1(new_n689), .B2(G1), .ZN(G364));
  INV_X1    g0490(.A(new_n652), .ZN(new_n691));
  INV_X1    g0491(.A(G13), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G20), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n209), .B1(new_n693), .B2(G45), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n637), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(G330), .B2(new_n636), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n233), .A2(new_n280), .ZN(new_n699));
  INV_X1    g0499(.A(G355), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(G116), .B2(new_n233), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n248), .A2(new_n307), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n233), .A2(new_n278), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n307), .B2(new_n229), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n701), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(G13), .A2(G33), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G20), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n230), .B1(G20), .B2(new_n340), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n696), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n210), .A2(new_n406), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G200), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(new_n369), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n210), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n716), .A2(new_n202), .B1(new_n205), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G190), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n713), .A2(G190), .A3(new_n329), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n280), .B1(new_n721), .B2(new_n351), .C1(new_n294), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n210), .A2(G179), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n369), .A3(G200), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G190), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(G87), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n206), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n719), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n724), .A2(new_n720), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G159), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n714), .A2(G190), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n732), .A2(KEYINPUT32), .B1(new_n733), .B2(G68), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n729), .B(new_n734), .C1(KEYINPUT32), .C2(new_n732), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n726), .B(KEYINPUT93), .Z(new_n736));
  AOI21_X1  g0536(.A(new_n280), .B1(new_n736), .B2(G303), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT94), .ZN(new_n738));
  INV_X1    g0538(.A(G326), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n716), .A2(new_n739), .B1(new_n740), .B2(new_n718), .ZN(new_n741));
  INV_X1    g0541(.A(new_n733), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT33), .B(G317), .Z(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n742), .A2(new_n743), .B1(new_n725), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n721), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G311), .A2(new_n747), .B1(new_n731), .B2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G322), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n746), .B(new_n748), .C1(new_n749), .C2(new_n722), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n738), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n712), .B1(new_n751), .B2(new_n709), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n708), .B(KEYINPUT95), .Z(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n636), .B2(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n698), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(G396));
  NOR2_X1   g0556(.A1(new_n709), .A2(new_n706), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n696), .B1(G77), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n722), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G143), .B1(new_n747), .B2(G159), .ZN(new_n761));
  INV_X1    g0561(.A(G137), .ZN(new_n762));
  INV_X1    g0562(.A(G150), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n761), .B1(new_n716), .B2(new_n762), .C1(new_n763), .C2(new_n742), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT96), .Z(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT34), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT34), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n278), .B1(new_n731), .B2(G132), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n768), .B1(new_n216), .B2(new_n725), .C1(new_n294), .C2(new_n718), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(G50), .B2(new_n736), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n736), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n206), .ZN(new_n773));
  INV_X1    g0573(.A(new_n718), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G97), .A2(new_n774), .B1(new_n715), .B2(G303), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n280), .B1(new_n747), .B2(G116), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n760), .A2(G294), .B1(new_n731), .B2(G311), .ZN(new_n777));
  INV_X1    g0577(.A(new_n725), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n733), .A2(G283), .B1(new_n778), .B2(G87), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n771), .B1(new_n773), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n759), .B1(new_n781), .B2(new_n709), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n424), .A2(new_n634), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n440), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n605), .B2(new_n783), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n782), .B1(new_n785), .B2(new_n707), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n626), .A2(new_n785), .A3(new_n643), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT97), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n785), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(new_n627), .B2(new_n634), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n687), .ZN(new_n793));
  INV_X1    g0593(.A(new_n696), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n792), .A2(new_n687), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n786), .B1(new_n795), .B2(new_n796), .ZN(G384));
  NOR2_X1   g0597(.A1(new_n693), .A2(new_n209), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n685), .B1(new_n596), .B2(new_n634), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n414), .A2(new_n415), .ZN(new_n800));
  INV_X1    g0600(.A(new_n401), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n415), .A2(new_n634), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n415), .B(new_n634), .C1(new_n414), .C2(new_n401), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n799), .A2(new_n805), .A3(new_n785), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(KEYINPUT40), .ZN(new_n807));
  AOI21_X1  g0607(.A(G200), .B1(new_n325), .B2(new_n327), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n288), .B(new_n304), .C1(new_n808), .C2(new_n324), .ZN(new_n809));
  INV_X1    g0609(.A(new_n304), .ZN(new_n810));
  INV_X1    g0610(.A(new_n285), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n279), .A2(new_n281), .ZN(new_n812));
  INV_X1    g0612(.A(new_n283), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n216), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n262), .A2(new_n274), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n276), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n287), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n811), .B1(new_n817), .B2(KEYINPUT101), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n284), .A2(new_n262), .A3(new_n274), .ZN(new_n819));
  AOI211_X1 g0619(.A(KEYINPUT101), .B(new_n301), .C1(new_n819), .C2(new_n276), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n810), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n341), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n809), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n632), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT37), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n305), .A2(new_n341), .ZN(new_n827));
  INV_X1    g0627(.A(new_n632), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n305), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT37), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .A4(new_n809), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n331), .A2(new_n336), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT80), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT80), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n600), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n825), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n838), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n301), .B1(new_n819), .B2(new_n276), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n285), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n304), .B1(new_n843), .B2(new_n820), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n828), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n608), .B2(new_n600), .ZN(new_n846));
  INV_X1    g0646(.A(new_n831), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n341), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n848), .A3(new_n809), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n849), .B2(KEYINPUT37), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n826), .A2(new_n831), .B1(new_n837), .B2(new_n825), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT102), .B1(new_n853), .B2(KEYINPUT38), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n807), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n827), .A2(new_n809), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n830), .A4(new_n829), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n827), .A2(new_n829), .A3(new_n809), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n831), .A2(KEYINPUT103), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n305), .B(new_n828), .C1(new_n345), .C2(new_n833), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(KEYINPUT38), .B2(new_n853), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT40), .B1(new_n865), .B2(new_n806), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n855), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n441), .A2(new_n799), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT105), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n671), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n869), .B2(new_n867), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT106), .Z(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  INV_X1    g0674(.A(new_n809), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n844), .B2(new_n341), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n830), .B1(new_n876), .B2(new_n845), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n347), .A2(new_n845), .B1(new_n877), .B2(new_n847), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n874), .B1(new_n878), .B2(new_n840), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n851), .A3(new_n839), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n601), .A2(new_n634), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n787), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n805), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n880), .A2(new_n885), .B1(new_n345), .B2(new_n632), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n880), .A2(KEYINPUT39), .B1(new_n865), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n414), .A2(new_n415), .A3(new_n643), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n441), .B1(new_n668), .B2(new_n669), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n612), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n798), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n873), .B2(new_n893), .ZN(new_n895));
  INV_X1    g0695(.A(new_n449), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(KEYINPUT35), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n897), .A2(G116), .A3(new_n231), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n229), .A2(G77), .A3(new_n257), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n903), .A2(KEYINPUT99), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n202), .A2(G68), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT100), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n692), .A2(G1), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n895), .B(new_n901), .C1(new_n908), .C2(new_n909), .ZN(G367));
  INV_X1    g0710(.A(new_n709), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n495), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n736), .A2(G116), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(KEYINPUT46), .ZN(new_n914));
  AOI22_X1  g0714(.A1(G107), .A2(new_n774), .B1(new_n715), .B2(G311), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n733), .A2(G294), .B1(new_n778), .B2(G97), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n280), .B1(new_n747), .B2(G283), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT111), .B(G317), .Z(new_n918));
  AOI22_X1  g0718(.A1(new_n760), .A2(G303), .B1(new_n731), .B2(new_n918), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n726), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n733), .A2(G159), .B1(new_n921), .B2(new_n272), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n216), .B2(new_n718), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n715), .A2(G143), .B1(new_n778), .B2(G77), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n760), .A2(G150), .B1(new_n747), .B2(G50), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n278), .B1(new_n731), .B2(G137), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n914), .A2(new_n920), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT47), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n911), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n710), .B1(new_n233), .B2(new_n420), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n244), .A2(new_n703), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n696), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT112), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n492), .A2(new_n643), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n517), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n563), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(new_n753), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n460), .A2(new_n643), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n614), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n482), .A2(new_n514), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(KEYINPUT107), .C1(new_n948), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n648), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  INV_X1    g0752(.A(new_n941), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n952), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n950), .A2(new_n650), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT42), .Z(new_n958));
  NAND3_X1  g0758(.A1(new_n947), .A2(new_n949), .A3(new_n623), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n634), .B1(new_n959), .B2(new_n514), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n955), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n650), .A2(new_n639), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n950), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT44), .B1(new_n963), .B2(new_n950), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n963), .A2(KEYINPUT44), .A3(new_n950), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n965), .A2(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n637), .A3(new_n647), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n648), .B1(new_n968), .B2(new_n967), .C1(new_n965), .C2(new_n966), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n636), .A2(G330), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT109), .ZN(new_n974));
  INV_X1    g0774(.A(new_n649), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n646), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n973), .B(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n650), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n689), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n689), .B1(new_n972), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n652), .B(KEYINPUT41), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n695), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n944), .B1(new_n962), .B2(new_n983), .ZN(G387));
  OAI21_X1  g0784(.A(new_n278), .B1(new_n730), .B2(new_n739), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n760), .A2(new_n918), .B1(new_n747), .B2(G303), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n733), .A2(G311), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n749), .C2(new_n716), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT48), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n718), .A2(new_n744), .B1(new_n726), .B2(new_n740), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT49), .Z(new_n995));
  AOI211_X1 g0795(.A(new_n985), .B(new_n995), .C1(G116), .C2(new_n778), .ZN(new_n996));
  INV_X1    g0796(.A(new_n420), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n774), .A2(new_n997), .B1(new_n778), .B2(G97), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n715), .A2(G159), .B1(new_n921), .B2(G77), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n760), .A2(G50), .B1(new_n747), .B2(G68), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n278), .B1(new_n731), .B2(G150), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n297), .A2(new_n742), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n709), .B1(new_n996), .B2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n699), .A2(new_n653), .B1(G107), .B2(new_n233), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n241), .A2(G45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n653), .ZN(new_n1009));
  AOI211_X1 g0809(.A(G45), .B(new_n1009), .C1(G68), .C2(G77), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n417), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n703), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1006), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1005), .B(new_n696), .C1(new_n711), .C2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n646), .B2(new_n942), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n978), .B2(new_n695), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n979), .A2(new_n691), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n978), .A2(new_n689), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(G393));
  OR2_X1    g0820(.A1(new_n972), .A2(new_n979), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n972), .A2(new_n979), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n691), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n278), .B1(new_n731), .B2(G143), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n216), .B2(new_n726), .C1(new_n727), .C2(new_n725), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT115), .Z(new_n1026));
  AOI22_X1  g0826(.A1(G150), .A2(new_n715), .B1(new_n760), .B2(G159), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT51), .Z(new_n1028));
  OAI22_X1  g0828(.A1(new_n718), .A2(new_n351), .B1(new_n721), .B2(new_n417), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G50), .B2(new_n733), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G317), .A2(new_n715), .B1(new_n760), .B2(G311), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT52), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n278), .B1(new_n730), .B2(new_n749), .C1(new_n721), .C2(new_n740), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n742), .A2(new_n579), .B1(new_n206), .B2(new_n725), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n718), .A2(new_n495), .B1(new_n726), .B2(new_n744), .ZN(new_n1036));
  OR4_X1    g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(KEYINPUT116), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT116), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n709), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n251), .A2(new_n703), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n710), .B1(new_n205), .B2(new_n233), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n696), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n950), .B2(new_n708), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n972), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n695), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1023), .A2(new_n1048), .ZN(G390));
  AOI21_X1  g0849(.A(new_n794), .B1(new_n297), .B2(new_n757), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n760), .A2(G116), .B1(new_n731), .B2(G294), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n278), .C1(new_n205), .C2(new_n721), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n774), .A2(G77), .B1(new_n778), .B2(G68), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n206), .B2(new_n742), .C1(new_n744), .C2(new_n716), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(G87), .C2(new_n736), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT54), .B(G143), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n774), .A2(G159), .B1(new_n747), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n762), .B2(new_n742), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT119), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n921), .A2(G150), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT53), .ZN(new_n1062));
  INV_X1    g0862(.A(G125), .ZN(new_n1063));
  INV_X1    g0863(.A(G132), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n280), .B1(new_n730), .B2(new_n1063), .C1(new_n722), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(G128), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n716), .A2(new_n1066), .B1(new_n202), .B2(new_n725), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1062), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1055), .B1(new_n1060), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1050), .B1(new_n1069), .B2(new_n911), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT120), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n707), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n888), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT39), .B1(new_n852), .B2(new_n854), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n865), .A2(new_n887), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n884), .A2(new_n889), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n846), .A2(new_n850), .A3(new_n840), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n634), .B1(new_n661), .B2(new_n666), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n881), .B1(new_n1079), .B2(new_n785), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n805), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n889), .B1(new_n1078), .B2(new_n864), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1077), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n799), .A2(G330), .A3(new_n785), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n686), .A2(new_n785), .A3(new_n805), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1077), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1073), .B1(new_n1090), .B2(new_n695), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n441), .A2(new_n686), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n891), .A2(new_n612), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1084), .A2(new_n1081), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1087), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n883), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1095), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT117), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n652), .B1(new_n1101), .B2(new_n1089), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1086), .A2(new_n1088), .A3(new_n1099), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1092), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1094), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT117), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1099), .A2(KEYINPUT117), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1077), .A2(new_n1087), .A3(new_n1082), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1087), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1108), .B(new_n1109), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  AND4_X1   g0912(.A1(new_n1092), .A2(new_n1112), .A3(new_n691), .A4(new_n1103), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1091), .B1(new_n1104), .B2(new_n1113), .ZN(G378));
  INV_X1    g0914(.A(new_n377), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n366), .A2(new_n632), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n377), .B1(new_n366), .B2(new_n632), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1072), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n696), .B1(G50), .B2(new_n758), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n280), .B(new_n469), .C1(new_n731), .C2(G283), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n774), .A2(G68), .B1(new_n921), .B2(G77), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n760), .A2(G107), .B1(new_n747), .B2(new_n997), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n715), .A2(G116), .B1(new_n778), .B2(new_n272), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n205), .C2(new_n742), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT58), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n202), .B1(G33), .B2(G41), .C1(new_n469), .C2(new_n280), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n742), .A2(new_n1064), .B1(new_n716), .B2(new_n1063), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n760), .A2(G128), .B1(new_n747), .B2(G137), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n726), .B2(new_n1056), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G150), .C2(new_n774), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT121), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n778), .A2(G159), .ZN(new_n1142));
  AOI211_X1 g0942(.A(G33), .B(G41), .C1(new_n731), .C2(G124), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1134), .B1(new_n1131), .B2(new_n1130), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1124), .B1(new_n1146), .B2(new_n709), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n671), .B(new_n1122), .C1(new_n855), .C2(new_n866), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1122), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n867), .B2(G330), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n890), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n889), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n852), .A2(new_n854), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1155), .A2(new_n884), .B1(new_n600), .B2(new_n828), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n799), .A2(new_n805), .A3(new_n785), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1078), .B2(new_n864), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n880), .A2(new_n807), .B1(new_n1159), .B2(KEYINPUT40), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1122), .B1(new_n1160), .B2(new_n671), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n867), .A2(G330), .A3(new_n1151), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1153), .A2(new_n1163), .A3(KEYINPUT122), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT122), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n890), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1149), .B1(new_n1167), .B2(new_n695), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT57), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1110), .A2(new_n1111), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT123), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1094), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT123), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1170), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n691), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1172), .B2(new_n1094), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1103), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1180), .B2(new_n1167), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1168), .B1(new_n1177), .B2(new_n1181), .ZN(G375));
  OAI211_X1 g0982(.A(new_n1101), .B(new_n982), .C1(new_n1106), .C2(new_n1105), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n694), .B(KEYINPUT124), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1081), .A2(new_n706), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n696), .B1(G68), .B2(new_n758), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n722), .A2(new_n762), .B1(new_n730), .B2(new_n1066), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n278), .B(new_n1187), .C1(G150), .C2(new_n747), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n736), .A2(G159), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n774), .A2(G50), .B1(new_n778), .B2(new_n272), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n715), .B1(new_n733), .B2(new_n1057), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n715), .A2(G294), .B1(new_n747), .B2(G107), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n495), .B2(new_n742), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n278), .B1(new_n730), .B2(new_n579), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G283), .B2(new_n760), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n774), .A2(new_n997), .B1(new_n778), .B2(G77), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n772), .C2(new_n205), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1192), .B1(new_n1195), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1186), .B1(new_n1200), .B2(new_n709), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1105), .A2(new_n1184), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1183), .A2(new_n1202), .ZN(G381));
  INV_X1    g1003(.A(G375), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1091), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1023), .A2(new_n1048), .ZN(new_n1208));
  INV_X1    g1008(.A(G384), .ZN(new_n1209));
  OR2_X1    g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(G387), .A3(G381), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1204), .A2(new_n1207), .A3(new_n1213), .ZN(G407));
  NAND2_X1  g1014(.A1(new_n633), .A2(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1204), .A2(new_n1207), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(G407), .A2(new_n1217), .A3(G213), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT126), .ZN(G409));
  AND2_X1   g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1211), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(G390), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1208), .B1(new_n1211), .B2(new_n1220), .ZN(new_n1223));
  INV_X1    g1023(.A(G387), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G378), .B(new_n1168), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1180), .A2(new_n1167), .A3(new_n982), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1153), .A2(new_n1163), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1149), .B1(new_n1232), .B2(new_n1184), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1207), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1215), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n652), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1239), .B2(new_n1238), .ZN(new_n1241));
  AOI21_X1  g1041(.A(G384), .B1(new_n1241), .B2(new_n1202), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(G384), .A3(new_n1202), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1216), .A2(G2897), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1245), .B(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1237), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1229), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1244), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(new_n1242), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1236), .A2(new_n1215), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT62), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1216), .B1(new_n1230), .B2(new_n1235), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT62), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1228), .B1(new_n1250), .B2(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1255), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT63), .B1(new_n1255), .B2(new_n1252), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1227), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT127), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1252), .B(new_n1246), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1249), .C1(new_n1264), .C2(new_n1255), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1259), .A2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1207), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1269), .A2(new_n1230), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1245), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1270), .A2(new_n1245), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1228), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1227), .A3(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(G402));
endmodule


