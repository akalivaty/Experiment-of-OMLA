//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1237, new_n1238, new_n1239;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  NOR2_X1   g0013(.A1(G257), .A2(G264), .ZN(new_n214));
  NOR3_X1   g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G20), .ZN(new_n220));
  INV_X1    g0020(.A(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n216), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G68), .A2(G238), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G50), .A2(G226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n229));
  INV_X1    g0029(.A(G116), .ZN(new_n230));
  INV_X1    g0030(.A(G270), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n228), .B(new_n232), .C1(G97), .C2(G257), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(G1), .B2(G20), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT66), .B(KEYINPUT1), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n224), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G87), .B(G97), .Z(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n256), .A2(new_n258), .B1(G20), .B2(new_n203), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n218), .ZN(new_n265));
  INV_X1    g0065(.A(G20), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n209), .A2(new_n266), .A3(G1), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(new_n265), .B1(new_n202), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n265), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n268), .B1(new_n202), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT9), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1698), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n278), .A2(G223), .B1(G222), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G77), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n275), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n287), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G226), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(G200), .B1(new_n297), .B2(KEYINPUT10), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n288), .A2(new_n292), .A3(new_n295), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT72), .B1(new_n299), .B2(G190), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT72), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n296), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n274), .B(new_n298), .C1(new_n300), .C2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n279), .A2(new_n281), .A3(G232), .A4(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n275), .A2(new_n309), .A3(G232), .A4(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n275), .A2(G226), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n287), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n294), .A2(G238), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n292), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT13), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n291), .B1(new_n314), .B2(new_n287), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n316), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(KEYINPUT75), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(new_n323), .A3(new_n320), .A4(new_n316), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(G200), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n258), .A2(G77), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n202), .B2(new_n262), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n266), .A2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n265), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  INV_X1    g0130(.A(G68), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(new_n272), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n209), .A2(G1), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n328), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT12), .Z(new_n336));
  NOR3_X1   g0136(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n318), .A2(G190), .A3(new_n321), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n325), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n322), .A2(G169), .A3(new_n324), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n318), .A2(G179), .A3(new_n321), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n322), .A2(new_n344), .A3(G169), .A4(new_n324), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n337), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n299), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n273), .C1(G169), .C2(new_n299), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n278), .A2(G238), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n282), .A2(G107), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n283), .A2(G232), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n291), .B1(new_n355), .B2(new_n287), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n294), .A2(G244), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n349), .A3(new_n357), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT15), .B(G87), .Z(new_n363));
  AOI22_X1  g0163(.A1(new_n256), .A2(new_n261), .B1(new_n363), .B2(new_n258), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n266), .B2(new_n285), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n265), .B1(new_n285), .B2(new_n267), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n272), .A2(new_n285), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT70), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT71), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n306), .A2(new_n348), .A3(new_n351), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  XNOR2_X1  g0174(.A(G58), .B(G68), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(G20), .B1(G159), .B2(new_n261), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT77), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n266), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT76), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n279), .A2(new_n281), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n279), .B2(new_n281), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n266), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n378), .B1(new_n386), .B2(new_n331), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n280), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT76), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n279), .A2(new_n281), .A3(new_n381), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n392), .B2(new_n266), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT77), .B(G68), .C1(new_n393), .C2(new_n380), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n374), .B(new_n377), .C1(new_n387), .C2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n385), .B1(new_n275), .B2(G20), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n396), .A2(new_n379), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n376), .B1(new_n397), .B2(new_n331), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n269), .B1(new_n398), .B2(new_n374), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT78), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n256), .A2(new_n271), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT79), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n267), .A2(new_n265), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n404), .B1(new_n267), .B2(new_n255), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n387), .A2(new_n394), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n376), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT78), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n399), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n401), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n275), .A2(G226), .A3(G1698), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(KEYINPUT80), .B1(G33), .B2(G87), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n283), .A2(G223), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(KEYINPUT80), .C2(new_n411), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT81), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n414), .A2(new_n415), .A3(new_n287), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n414), .B2(new_n287), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n291), .B1(new_n294), .B2(G232), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n349), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n287), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n419), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n418), .A2(new_n420), .B1(new_n359), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n410), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n410), .A2(KEYINPUT18), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OR2_X1    g0228(.A1(KEYINPUT82), .A2(G190), .ZN(new_n429));
  NAND2_X1  g0229(.A1(KEYINPUT82), .A2(G190), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n419), .B(new_n431), .C1(new_n416), .C2(new_n417), .ZN(new_n432));
  INV_X1    g0232(.A(G200), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n401), .A2(new_n435), .A3(new_n405), .A4(new_n409), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT17), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n356), .B2(new_n357), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n370), .B1(new_n302), .B2(new_n358), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n428), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n373), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n275), .A2(new_n266), .A3(G68), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT86), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT19), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(new_n266), .A3(G33), .A4(G97), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G87), .A2(G97), .ZN(new_n447));
  INV_X1    g0247(.A(G107), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n447), .A2(new_n448), .B1(new_n313), .B2(new_n266), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n449), .B2(new_n445), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n275), .A2(KEYINPUT86), .A3(new_n266), .A4(G68), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n265), .ZN(new_n453));
  INV_X1    g0253(.A(new_n363), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n267), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n404), .B1(G1), .B2(new_n257), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G87), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n453), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(new_n290), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n293), .A2(G250), .A3(new_n462), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n283), .A2(G238), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n279), .A2(new_n281), .A3(G244), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT85), .B1(new_n467), .B2(new_n311), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT85), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n275), .A2(new_n469), .A3(G244), .A4(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  AOI211_X1 g0272(.A(new_n463), .B(new_n465), .C1(new_n472), .C2(new_n287), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n459), .B1(new_n473), .B2(new_n433), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT87), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT87), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n459), .B(new_n476), .C1(new_n473), .C2(new_n433), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(G190), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n448), .A2(G20), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT23), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n275), .A2(new_n266), .A3(G87), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(KEYINPUT91), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n484), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n275), .A2(new_n486), .A3(new_n266), .A4(G87), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n481), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n258), .A2(G116), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n265), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n480), .A2(G1), .A3(new_n209), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT25), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n457), .A2(G107), .B1(new_n495), .B2(new_n494), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G257), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G1698), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n275), .B(new_n500), .C1(G250), .C2(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G294), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n287), .ZN(new_n504));
  AND2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  NOR2_X1   g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n461), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n293), .A2(G264), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g0310(.A1(new_n507), .A2(new_n290), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT92), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n293), .B1(new_n501), .B2(new_n502), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n504), .A2(new_n509), .A3(new_n511), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n515), .A2(new_n349), .B1(new_n516), .B2(new_n359), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n498), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n473), .A2(new_n349), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n453), .B(new_n455), .C1(new_n454), .C2(new_n456), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(G169), .C2(new_n473), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n479), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n267), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n456), .A2(new_n523), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n448), .B1(new_n396), .B2(new_n379), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n523), .A2(new_n448), .ZN(new_n530));
  NOR2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n448), .A2(KEYINPUT6), .A3(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n266), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n262), .A2(new_n285), .ZN(new_n535));
  OR3_X1    g0335(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n527), .B1(new_n536), .B2(new_n265), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n528), .A2(new_n534), .A3(new_n535), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n538), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n524), .B(new_n526), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT4), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n467), .A2(new_n541), .B1(G33), .B2(G283), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n275), .A2(KEYINPUT4), .A3(G244), .A4(new_n311), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n275), .B2(G250), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n311), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n287), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n293), .A2(new_n507), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G257), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n546), .A2(G190), .A3(new_n511), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT84), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n545), .A2(new_n287), .B1(G257), .B2(new_n547), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(G190), .A4(new_n511), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n546), .A2(new_n511), .A3(new_n548), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n433), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n540), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n546), .A2(new_n511), .A3(new_n548), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n359), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n551), .A2(new_n349), .A3(new_n511), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n524), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n536), .A2(new_n527), .A3(new_n265), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT83), .B1(new_n538), .B2(new_n269), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n526), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n515), .A2(new_n433), .B1(new_n516), .B2(new_n302), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n498), .A2(new_n567), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n557), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n266), .C1(G33), .C2(new_n523), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(new_n265), .C1(new_n266), .C2(G116), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT88), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n577), .A3(new_n573), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n334), .A2(G20), .A3(new_n230), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n457), .A2(G116), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G303), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n282), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G264), .A2(G1698), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n499), .B2(G1698), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n287), .C1(new_n282), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n293), .A2(new_n507), .A3(G270), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n511), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G200), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n590), .A2(new_n431), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n583), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT90), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n590), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(new_n359), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n582), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT89), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n582), .A2(new_n597), .A3(KEYINPUT89), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n596), .A2(G179), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n596), .A2(new_n601), .A3(new_n359), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n582), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n595), .A2(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n441), .A2(new_n522), .A3(new_n569), .A4(new_n609), .ZN(G372));
  NAND3_X1  g0410(.A1(new_n479), .A2(new_n566), .A3(new_n521), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT26), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(new_n518), .A3(new_n607), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n498), .A2(new_n567), .ZN(new_n614));
  INV_X1    g0414(.A(new_n566), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n562), .B(new_n525), .C1(new_n563), .C2(new_n564), .ZN(new_n616));
  INV_X1    g0416(.A(new_n556), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n550), .A4(new_n553), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n478), .B(new_n459), .C1(new_n433), .C2(new_n473), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n521), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n612), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n621), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT93), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(new_n616), .B2(new_n561), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n540), .A2(KEYINPUT93), .A3(new_n560), .A4(new_n559), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n521), .B1(new_n627), .B2(KEYINPUT26), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n441), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n351), .ZN(new_n631));
  INV_X1    g0431(.A(new_n372), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n339), .B1(new_n347), .B2(new_n346), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n401), .A2(new_n409), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT17), .A3(new_n435), .A4(new_n405), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT17), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n436), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n428), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n631), .B1(new_n639), .B2(new_n306), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n640), .ZN(G369));
  NAND3_X1  g0441(.A1(new_n270), .A2(new_n266), .A3(G13), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n582), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n608), .B(new_n609), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n647), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n498), .A2(new_n517), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n498), .A2(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n614), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n518), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n647), .B1(new_n603), .B2(new_n607), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n654), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(G399));
  NOR2_X1   g0461(.A1(new_n212), .A2(G41), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n447), .A2(new_n448), .A3(new_n230), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n222), .B2(new_n663), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n569), .A2(new_n623), .A3(new_n613), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n627), .A2(KEYINPUT26), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n611), .A2(KEYINPUT26), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n521), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n652), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT29), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n629), .A2(new_n652), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(KEYINPUT29), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n609), .A2(new_n569), .A3(new_n522), .A4(new_n652), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n510), .A2(new_n514), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n678), .A2(new_n605), .A3(new_n555), .A4(new_n473), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT30), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n555), .A2(new_n473), .A3(G179), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n515), .A3(new_n590), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(KEYINPUT30), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n647), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(KEYINPUT31), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n676), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n668), .B1(new_n689), .B2(G1), .ZN(G364));
  OR2_X1    g0490(.A1(new_n649), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n266), .A2(G13), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT94), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n270), .B1(new_n694), .B2(G45), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n662), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n691), .A2(new_n650), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G179), .A2(G200), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n266), .B1(new_n700), .B2(G190), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G97), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(G20), .A3(new_n302), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G159), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n266), .A2(new_n349), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G200), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G190), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI221_X1 g0510(.A(new_n703), .B1(new_n706), .B2(KEYINPUT32), .C1(new_n710), .C2(new_n331), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n708), .A2(new_n431), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G50), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n302), .A3(new_n433), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n433), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n431), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G58), .ZN(new_n718));
  OAI221_X1 g0518(.A(new_n713), .B1(new_n285), .B2(new_n714), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n711), .B(new_n719), .C1(KEYINPUT32), .C2(new_n706), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n433), .A2(G179), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(G20), .A3(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G87), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(G20), .A3(new_n302), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT98), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT98), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT99), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G107), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n720), .A2(new_n275), .A3(new_n724), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(G317), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n733), .A2(new_n709), .B1(G322), .B2(new_n716), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT101), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n275), .B1(new_n705), .B2(G329), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n584), .B2(new_n722), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  INV_X1    g0538(.A(G294), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n714), .A2(new_n738), .B1(new_n701), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n729), .ZN(new_n742));
  INV_X1    g0542(.A(G283), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n735), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n712), .A2(G326), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n731), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n218), .B1(G20), .B2(new_n359), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n209), .A2(new_n257), .A3(KEYINPUT96), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT96), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G13), .B2(G33), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n748), .B1(new_n649), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n392), .A2(new_n211), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n221), .A2(new_n460), .A3(G50), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(new_n460), .C2(new_n250), .ZN(new_n760));
  INV_X1    g0560(.A(G355), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n211), .A2(new_n275), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n760), .B1(G116), .B2(new_n211), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n754), .A2(new_n747), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n698), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  OAI21_X1  g0566(.A(new_n699), .B1(new_n756), .B2(new_n766), .ZN(G396));
  AND4_X1   g0567(.A1(new_n371), .A2(new_n360), .A3(new_n361), .A4(new_n652), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n439), .A2(new_n438), .B1(new_n370), .B2(new_n652), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(new_n769), .B2(new_n372), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n770), .B(KEYINPUT104), .ZN(new_n772));
  MUX2_X1   g0572(.A(new_n771), .B(new_n772), .S(new_n675), .Z(new_n773));
  INV_X1    g0573(.A(new_n688), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n698), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n282), .B1(new_n704), .B2(new_n738), .C1(new_n722), .C2(new_n448), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n710), .A2(new_n743), .B1(new_n714), .B2(new_n230), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n729), .C2(G87), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n703), .B1(new_n717), .B2(new_n739), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT102), .ZN(new_n781));
  INV_X1    g0581(.A(new_n712), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n779), .B(new_n781), .C1(new_n584), .C2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT103), .Z(new_n784));
  INV_X1    g0584(.A(new_n392), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n202), .B2(new_n722), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n742), .A2(new_n331), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G58), .C2(new_n702), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G143), .A2(new_n716), .B1(new_n709), .B2(G150), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n782), .C1(new_n791), .C2(new_n714), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT34), .ZN(new_n793));
  INV_X1    g0593(.A(G132), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n788), .B(new_n793), .C1(new_n794), .C2(new_n704), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n698), .B1(new_n796), .B2(new_n747), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n752), .A2(new_n747), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n797), .B1(G77), .B2(new_n799), .C1(new_n753), .C2(new_n770), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n776), .A2(new_n800), .ZN(G384));
  INV_X1    g0601(.A(new_n645), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n410), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n424), .A2(new_n803), .A3(new_n436), .ZN(new_n804));
  XOR2_X1   g0604(.A(KEYINPUT107), .B(KEYINPUT37), .Z(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT108), .ZN(new_n807));
  INV_X1    g0607(.A(new_n805), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n424), .A2(new_n803), .A3(new_n436), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n803), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n410), .A2(KEYINPUT18), .A3(new_n423), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT18), .B1(new_n410), .B2(new_n423), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n814), .B2(new_n638), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n809), .A2(new_n807), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n810), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n377), .B1(new_n387), .B2(new_n394), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n265), .B1(new_n820), .B2(KEYINPUT16), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n405), .B1(new_n821), .B2(new_n395), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n802), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n814), .B2(new_n638), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n423), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(new_n823), .A3(new_n436), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n809), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n825), .A2(KEYINPUT38), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT109), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n637), .B(new_n635), .C1(new_n812), .C2(new_n813), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(new_n824), .B1(new_n809), .B2(new_n828), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT109), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT38), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n819), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n346), .A2(new_n347), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n647), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n823), .B1(new_n428), .B2(new_n437), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n828), .A2(new_n809), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n818), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n843), .A2(KEYINPUT39), .A3(new_n830), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT106), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n347), .A2(new_n647), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n348), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n348), .B2(new_n847), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n652), .B(new_n770), .C1(new_n622), .C2(new_n628), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT105), .ZN(new_n853));
  INV_X1    g0653(.A(new_n768), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n851), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n830), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n814), .A2(new_n645), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n846), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n676), .A2(new_n441), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n640), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n864), .B(new_n866), .Z(new_n867));
  OAI21_X1  g0667(.A(new_n770), .B1(new_n849), .B2(new_n850), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n686), .A2(new_n687), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n858), .B2(new_n859), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n873), .A2(KEYINPUT110), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(KEYINPUT110), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n373), .A2(new_n440), .A3(new_n869), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G330), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n867), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n270), .B2(new_n694), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n532), .A2(new_n533), .ZN(new_n883));
  OAI211_X1 g0683(.A(G20), .B(new_n219), .C1(new_n883), .C2(KEYINPUT35), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n230), .B(new_n884), .C1(KEYINPUT35), .C2(new_n883), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  OAI21_X1  g0686(.A(G77), .B1(new_n718), .B2(new_n331), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n222), .A2(new_n887), .B1(G50), .B2(new_n331), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(G1), .A3(new_n209), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n882), .A2(new_n886), .A3(new_n889), .ZN(G367));
  OAI22_X1  g0690(.A1(new_n714), .A2(new_n743), .B1(new_n701), .B2(new_n448), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n722), .A2(new_n230), .ZN(new_n894));
  AOI22_X1  g0694(.A1(KEYINPUT46), .A2(new_n894), .B1(new_n712), .B2(G311), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n785), .B1(G317), .B2(new_n705), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n584), .B2(new_n717), .ZN(new_n898));
  INV_X1    g0698(.A(new_n728), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(G97), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(KEYINPUT46), .B2(new_n894), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n896), .B(new_n901), .C1(G294), .C2(new_n709), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n705), .A2(G137), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n702), .A2(G68), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n904), .B1(new_n202), .B2(new_n714), .C1(new_n710), .C2(new_n791), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n282), .B1(new_n723), .B2(G58), .ZN(new_n906));
  INV_X1    g0706(.A(G143), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n906), .B1(new_n782), .B2(new_n907), .C1(new_n260), .C2(new_n717), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n905), .B(new_n908), .C1(G77), .C2(new_n899), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n902), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT47), .Z(new_n911));
  AOI21_X1  g0711(.A(new_n698), .B1(new_n911), .B2(new_n747), .ZN(new_n912));
  INV_X1    g0712(.A(new_n758), .ZN(new_n913));
  OAI221_X1 g0713(.A(new_n764), .B1(new_n211), .B2(new_n454), .C1(new_n913), .C2(new_n242), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n459), .A2(new_n652), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT111), .Z(new_n916));
  INV_X1    g0716(.A(new_n521), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n621), .B2(new_n916), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n912), .B(new_n914), .C1(new_n755), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n615), .B(new_n618), .C1(new_n616), .C2(new_n652), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n615), .B2(new_n652), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n660), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT45), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n660), .A2(new_n922), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n658), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n658), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n657), .B(new_n659), .Z(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(new_n650), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n689), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n689), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n662), .B(KEYINPUT41), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n696), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n928), .A2(new_n922), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n657), .A2(new_n659), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n921), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT42), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n615), .B1(new_n921), .B2(new_n518), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n652), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n928), .A2(new_n922), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n944), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n950), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n920), .B1(new_n937), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT113), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT113), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n920), .C1(new_n937), .C2(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(G387));
  NAND2_X1  g0758(.A1(new_n933), .A2(new_n696), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT114), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G311), .A2(new_n709), .B1(new_n716), .B2(G317), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n584), .B2(new_n714), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G322), .B2(new_n712), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT48), .Z(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n743), .B2(new_n701), .C1(new_n739), .C2(new_n722), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT49), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n705), .A2(G326), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n785), .B1(new_n899), .B2(G116), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n782), .A2(new_n791), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n710), .A2(new_n255), .B1(new_n714), .B2(new_n331), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n785), .B1(new_n260), .B2(new_n704), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G77), .C2(new_n723), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n716), .A2(G50), .B1(new_n363), .B2(new_n702), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT117), .Z(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n523), .C2(new_n742), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n971), .B1(new_n972), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n747), .ZN(new_n980));
  AOI211_X1 g0780(.A(G45), .B(new_n664), .C1(G68), .C2(G77), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT50), .B1(new_n255), .B2(G50), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(KEYINPUT115), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n255), .A2(KEYINPUT50), .A3(G50), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n758), .C1(new_n460), .C2(new_n246), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(G107), .B2(new_n211), .C1(new_n665), .C2(new_n762), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n698), .B1(new_n989), .B2(new_n764), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT116), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n980), .B(new_n991), .C1(new_n657), .C2(new_n755), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n934), .A2(new_n662), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT118), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n689), .A2(new_n933), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT119), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n996), .A2(new_n997), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n960), .B(new_n992), .C1(new_n999), .C2(new_n1000), .ZN(G393));
  AOI21_X1  g0801(.A(new_n663), .B1(new_n931), .B2(new_n934), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n931), .B2(new_n934), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n764), .B1(new_n523), .B2(new_n211), .C1(new_n913), .C2(new_n253), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G311), .A2(new_n716), .B1(new_n712), .B2(G317), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT52), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n709), .A2(G303), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n282), .B1(new_n722), .B2(new_n743), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n714), .A2(new_n739), .B1(new_n701), .B2(new_n230), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(G322), .C2(new_n705), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1006), .A2(new_n730), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n729), .A2(G87), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n785), .B1(new_n907), .B2(new_n704), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT121), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n710), .A2(new_n202), .B1(new_n714), .B2(new_n255), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1012), .B(new_n1016), .C1(new_n331), .C2(new_n722), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G150), .A2(new_n712), .B1(new_n716), .B2(G159), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n702), .A2(G77), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n698), .B1(new_n1023), .B2(new_n747), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1004), .B(new_n1024), .C1(new_n922), .C2(new_n755), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1003), .B(new_n1025), .C1(new_n695), .C2(new_n931), .ZN(G390));
  NAND2_X1  g0826(.A1(new_n769), .A2(new_n372), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n854), .B1(new_n673), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n840), .B1(new_n1029), .B2(new_n851), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n836), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n844), .B1(new_n836), .B2(new_n837), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n852), .A2(new_n854), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT105), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n840), .B1(new_n1036), .B2(new_n851), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1031), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n688), .A2(new_n770), .A3(new_n851), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1031), .B(new_n1039), .C1(new_n1032), .C2(new_n1037), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n878), .A2(G330), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n640), .A3(new_n865), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n851), .B1(new_n688), .B2(new_n772), .ZN(new_n1045));
  OR3_X1    g0845(.A1(new_n1040), .A2(new_n1029), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n851), .B1(new_n688), .B2(new_n770), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1036), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1044), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1041), .A2(new_n1042), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT122), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1041), .A2(new_n1049), .A3(KEYINPUT122), .A4(new_n1042), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n857), .B1(new_n839), .B2(new_n647), .ZN(new_n1055));
  AND4_X1   g0855(.A1(new_n834), .A2(new_n825), .A3(KEYINPUT38), .A4(new_n829), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n834), .B1(new_n833), .B2(KEYINPUT38), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT39), .B1(new_n1058), .B2(new_n819), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1055), .B1(new_n1059), .B2(new_n844), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1039), .B1(new_n1060), .B2(new_n1031), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1042), .ZN(new_n1062));
  OAI21_X1  g0862(.A(KEYINPUT123), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1049), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT123), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1041), .A2(new_n1065), .A3(new_n1042), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1054), .A2(new_n1067), .A3(new_n662), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G107), .A2(new_n709), .B1(new_n716), .B2(G116), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n724), .C1(new_n523), .C2(new_n714), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1021), .B1(new_n739), .B2(new_n704), .C1(new_n782), .C2(new_n743), .ZN(new_n1071));
  OR4_X1    g0871(.A1(new_n275), .A2(new_n787), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT54), .B(G143), .Z(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n714), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n723), .A2(G150), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT53), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1075), .B(new_n1077), .C1(G137), .C2(new_n709), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n705), .A2(G125), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n899), .A2(G50), .ZN(new_n1080));
  INV_X1    g0880(.A(G128), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n782), .A2(new_n1081), .B1(new_n791), .B2(new_n701), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n282), .B(new_n1082), .C1(G132), .C2(new_n716), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1072), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT124), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n698), .B1(new_n1086), .B2(new_n747), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n256), .B2(new_n799), .C1(new_n1032), .C2(new_n753), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n696), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1068), .A2(new_n1091), .ZN(G378));
  INV_X1    g0892(.A(new_n1044), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1054), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n306), .A2(new_n351), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT55), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n273), .A2(new_n802), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT56), .Z(new_n1098));
  XNOR2_X1  g0898(.A(new_n1096), .B(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n871), .A2(new_n876), .A3(G330), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n864), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n871), .A2(new_n876), .A3(G330), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n861), .B1(new_n1032), .B2(new_n840), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n863), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n864), .A2(new_n1101), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n863), .A3(new_n1103), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n1108), .A3(new_n1099), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1094), .A2(KEYINPUT57), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT57), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1044), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1107), .A2(new_n1099), .A3(new_n1108), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1099), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1111), .A2(new_n1117), .A3(new_n662), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1099), .A2(new_n752), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n798), .A2(new_n202), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G107), .A2(new_n716), .B1(new_n712), .B2(G116), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1121), .B1(new_n523), .B2(new_n710), .C1(new_n454), .C2(new_n714), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n728), .A2(new_n718), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n392), .B(new_n904), .C1(new_n743), .C2(new_n704), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1123), .A2(G41), .A3(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1122), .B(new_n1125), .C1(G77), .C2(new_n723), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT58), .Z(new_n1127));
  OAI22_X1  g0927(.A1(new_n1074), .A2(new_n722), .B1(new_n714), .B2(new_n790), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G125), .A2(new_n712), .B1(new_n709), .B2(G132), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1081), .B2(new_n717), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G150), .C2(new_n702), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT59), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G41), .B1(new_n899), .B2(G159), .ZN(new_n1133));
  AOI21_X1  g0933(.A(G33), .B1(new_n705), .B2(G124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(G41), .B1(new_n785), .B2(G33), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1127), .B(new_n1135), .C1(G50), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n698), .B1(new_n1137), .B2(new_n747), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1119), .A2(new_n1120), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1110), .B2(new_n696), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1118), .A2(new_n1140), .ZN(G375));
  AND2_X1   g0941(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1044), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n936), .A3(new_n1064), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G137), .A2(new_n716), .B1(new_n709), .B2(new_n1073), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n794), .B2(new_n782), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT125), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n785), .B1(new_n791), .B2(new_n722), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n714), .A2(new_n260), .B1(new_n701), .B2(new_n202), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1123), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1147), .B(new_n1150), .C1(new_n1081), .C2(new_n704), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G283), .A2(new_n716), .B1(new_n712), .B2(G294), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n448), .B2(new_n714), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n710), .A2(new_n230), .B1(new_n454), .B2(new_n701), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n282), .B1(new_n704), .B2(new_n584), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n523), .B2(new_n722), .C1(new_n742), .C2(new_n285), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n747), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(G68), .B2(new_n799), .C1(new_n851), .C2(new_n753), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(new_n698), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1142), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n696), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1144), .A2(new_n1163), .ZN(G381));
  NOR4_X1   g0964(.A1(G387), .A2(G384), .A3(G390), .A4(G381), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(G393), .A2(G396), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1140), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1165), .A2(new_n1118), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT126), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(G407));
  NAND3_X1  g0970(.A1(new_n1140), .A2(new_n1068), .A3(new_n1091), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n663), .B1(new_n1172), .B2(KEYINPUT57), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1173), .B2(new_n1117), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n646), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1177));
  OAI211_X1 g0977(.A(G213), .B(new_n1175), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT127), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(G407), .A2(KEYINPUT127), .A3(G213), .A4(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(G409));
  XNOR2_X1  g0982(.A(G393), .B(G396), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n954), .A2(G390), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n954), .A2(G390), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(G387), .B2(G390), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1183), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT61), .ZN(new_n1193));
  INV_X1    g0993(.A(G378), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1118), .B2(new_n1140), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1094), .A2(new_n936), .A3(new_n1110), .ZN(new_n1196));
  INV_X1    g0996(.A(G213), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n1196), .A2(new_n1171), .B1(new_n1197), .B2(G343), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT60), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1143), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n1044), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n662), .A3(new_n1064), .A4(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G384), .B1(new_n1202), .B2(new_n1163), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(G384), .A3(new_n1163), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1195), .A2(new_n1198), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT62), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1193), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1197), .A2(G343), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(G2897), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1205), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1211), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1203), .A3(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1172), .A2(new_n936), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1210), .B1(new_n1167), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1206), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1140), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1173), .B2(new_n1117), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1219), .B(new_n1220), .C1(new_n1222), .C2(new_n1194), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT62), .B1(new_n1217), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1192), .B1(new_n1209), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1214), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1204), .A2(new_n1205), .A3(new_n1211), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G375), .A2(G378), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n1229), .B2(new_n1219), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT63), .B1(new_n1230), .B2(new_n1207), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1192), .A2(KEYINPUT61), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT63), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1223), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1225), .A2(new_n1235), .ZN(G405));
  OR3_X1    g1036(.A1(new_n1195), .A2(new_n1174), .A3(new_n1220), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1220), .B1(new_n1195), .B2(new_n1174), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(new_n1191), .ZN(G402));
endmodule


