//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(KEYINPUT2), .B2(G113), .ZN(new_n193));
  AOI22_X1  g007(.A1(new_n191), .A2(new_n193), .B1(KEYINPUT2), .B2(G113), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n194), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT0), .A4(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT0), .B(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G137), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(G134), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g034(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n212), .C2(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G131), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n219), .B1(new_n214), .B2(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n217), .A3(new_n219), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n216), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n211), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n213), .A2(new_n215), .ZN(new_n231));
  AOI211_X1 g045(.A(G131), .B(new_n231), .C1(new_n225), .C2(new_n226), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n233));
  OAI211_X1 g047(.A(G128), .B(new_n233), .C1(new_n207), .C2(new_n208), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n218), .A2(new_n215), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n203), .B(new_n205), .C1(KEYINPUT1), .C2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n234), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n201), .B1(new_n230), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n211), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n228), .B1(new_n227), .B2(new_n216), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n232), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n194), .B(new_n199), .ZN(new_n245));
  INV_X1    g059(.A(new_n239), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n229), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n188), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n223), .A2(new_n229), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n250), .A2(new_n242), .B1(new_n229), .B2(new_n246), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n251), .B2(new_n245), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT70), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n230), .A2(new_n240), .A3(new_n201), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n245), .B1(new_n244), .B2(new_n247), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT28), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n253), .A2(new_n258), .A3(KEYINPUT29), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n249), .A2(new_n252), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n267), .B2(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n248), .A2(new_n188), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n272), .B(new_n273), .C1(new_n230), .C2(new_n240), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n244), .A2(KEYINPUT65), .A3(new_n271), .A4(new_n247), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n245), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n266), .B1(new_n276), .B2(new_n254), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n187), .B(new_n264), .C1(new_n268), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G472), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT67), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n275), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n201), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n263), .A4(new_n248), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n266), .B1(new_n249), .B2(new_n252), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n276), .A2(new_n254), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n286), .B1(new_n290), .B2(new_n263), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT32), .B(new_n283), .C1(new_n289), .C2(new_n291), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n280), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(G217), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(G234), .ZN(new_n299));
  XOR2_X1   g113(.A(new_n299), .B(KEYINPUT71), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G125), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G140), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT16), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n308), .B1(new_n303), .B2(KEYINPUT16), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G146), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n305), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT76), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n202), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n195), .A2(G128), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT72), .A3(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n237), .A2(KEYINPUT73), .A3(G119), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n237), .A2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT72), .B1(new_n319), .B2(KEYINPUT23), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  OAI22_X1  g141(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(new_n322), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n322), .A2(new_n319), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  OAI22_X1  g144(.A1(new_n328), .A2(G110), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G137), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(KEYINPUT74), .A3(G110), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT74), .B1(new_n328), .B2(G110), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n202), .B(new_n306), .C1(new_n307), .C2(new_n309), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n311), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n329), .A2(new_n330), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n332), .B(new_n336), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n339), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n337), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n347), .A2(new_n348), .B1(new_n331), .B2(new_n318), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n336), .B(KEYINPUT77), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n345), .B(new_n187), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n332), .B1(new_n340), .B2(new_n344), .ZN(new_n354));
  INV_X1    g168(.A(new_n350), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(KEYINPUT25), .A3(new_n187), .A4(new_n345), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n301), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n345), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n301), .A2(new_n187), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n296), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT87), .A2(G143), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT87), .A2(G143), .ZN(new_n365));
  OAI211_X1 g179(.A(G214), .B(new_n259), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G237), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n334), .A3(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT87), .A2(G143), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n228), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT17), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n311), .A2(new_n341), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT89), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n311), .A2(new_n372), .A3(new_n375), .A4(new_n341), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n366), .A2(new_n228), .A3(new_n370), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n377), .A2(new_n371), .A3(KEYINPUT17), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n317), .B1(new_n202), .B2(new_n315), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n371), .A2(KEYINPUT18), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT18), .A2(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n366), .A2(new_n370), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(G113), .B(G122), .Z(new_n387));
  XOR2_X1   g201(.A(KEYINPUT88), .B(G104), .Z(new_n388));
  XOR2_X1   g202(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n312), .A2(KEYINPUT19), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n314), .A2(new_n316), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(KEYINPUT19), .ZN(new_n393));
  OAI221_X1 g207(.A(new_n311), .B1(new_n371), .B2(new_n377), .C1(new_n393), .C2(G146), .ZN(new_n394));
  INV_X1    g208(.A(new_n385), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n390), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n386), .A2(new_n390), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n397), .A2(KEYINPUT90), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT90), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n385), .A3(new_n389), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n378), .B1(new_n373), .B2(KEYINPUT89), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n395), .B1(new_n403), .B2(new_n376), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n399), .C1(new_n404), .C2(new_n389), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n401), .B1(new_n405), .B2(KEYINPUT20), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n404), .B2(new_n412), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G475), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT92), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n410), .A2(KEYINPUT92), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n204), .A2(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n237), .A2(G143), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n214), .ZN(new_n423));
  XNOR2_X1  g237(.A(G116), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(G107), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n424), .ZN(new_n428));
  OAI211_X1 g242(.A(G107), .B(new_n427), .C1(new_n428), .C2(KEYINPUT14), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n424), .B(new_n425), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n214), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n420), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n204), .A2(KEYINPUT13), .A3(G128), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(new_n421), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n431), .B(new_n432), .C1(new_n214), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n438), .A2(new_n298), .A3(G953), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n430), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n430), .B2(new_n437), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n187), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G478), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT15), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G952), .A3(new_n334), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(G898), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n418), .A2(new_n419), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G110), .B(G122), .ZN(new_n459));
  INV_X1    g273(.A(G104), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT3), .B1(new_n460), .B2(G107), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n425), .A3(G104), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(G107), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(G101), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(G101), .ZN(new_n468));
  INV_X1    g282(.A(G101), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n461), .A2(new_n463), .A3(new_n469), .A4(new_n464), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(KEYINPUT4), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n201), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G104), .B(G107), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT78), .B1(new_n473), .B2(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n425), .A2(G104), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n464), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT78), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(G101), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n194), .A2(new_n200), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT5), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(G113), .C1(KEYINPUT5), .C2(new_n196), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n470), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n459), .B1(new_n472), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT6), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n465), .A2(G101), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n467), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n483), .B(new_n459), .C1(new_n489), .C2(new_n245), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n472), .A2(new_n492), .A3(new_n459), .A4(new_n483), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n486), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n485), .B1(new_n494), .B2(new_n484), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n211), .A2(G125), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n234), .A2(new_n238), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n498), .B2(G125), .ZN(new_n499));
  INV_X1    g313(.A(G224), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n499), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT85), .Z(new_n505));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(new_n500), .B2(G953), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n499), .B(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n477), .B1(new_n476), .B2(G101), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT78), .B(new_n469), .C1(new_n475), .C2(new_n464), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n470), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n480), .A2(new_n482), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G113), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(KEYINPUT83), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n481), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(new_n480), .A3(new_n470), .A4(new_n479), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT84), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n459), .B(KEYINPUT8), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n507), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n491), .A2(new_n493), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n503), .A2(new_n505), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n505), .B1(new_n503), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(G214), .B1(G237), .B2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G469), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n510), .B2(new_n497), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n471), .A2(new_n242), .A3(new_n467), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n498), .A2(new_n479), .A3(KEYINPUT10), .A4(new_n470), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n250), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G140), .ZN(new_n540));
  INV_X1    g354(.A(G227), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(G953), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n540), .B(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT79), .B1(new_n232), .B2(new_n243), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT79), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n223), .A2(new_n546), .A3(new_n229), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n539), .B(new_n544), .C1(new_n538), .C2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n510), .A2(new_n497), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n479), .A2(new_n470), .B1(new_n238), .B2(new_n234), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n250), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT12), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT12), .B(new_n250), .C1(new_n550), .C2(new_n551), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n556));
  INV_X1    g370(.A(new_n548), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n549), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n533), .B1(new_n559), .B2(new_n187), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n544), .B1(new_n538), .B2(new_n548), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT81), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n554), .A2(new_n555), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT81), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n544), .C1(new_n538), .C2(new_n548), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n556), .A2(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n539), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n543), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT80), .B(G469), .Z(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n187), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n532), .B1(new_n561), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n530), .A2(new_n575), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n363), .A2(new_n458), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n469), .ZN(G3));
  OAI21_X1  g392(.A(new_n187), .B1(new_n289), .B2(new_n291), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  AND4_X1   g394(.A1(new_n292), .A2(new_n575), .A3(new_n362), .A4(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n440), .B2(new_n441), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT33), .Z(new_n584));
  NOR2_X1   g398(.A1(new_n444), .A2(G902), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n584), .A2(new_n585), .B1(new_n444), .B2(new_n442), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n418), .B2(new_n419), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n503), .A2(new_n525), .ZN(new_n588));
  INV_X1    g402(.A(new_n505), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n503), .A2(new_n505), .A3(new_n525), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n528), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n456), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n581), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n593), .ZN(new_n597));
  INV_X1    g411(.A(new_n449), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(G475), .B2(new_n414), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n405), .B(new_n408), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT35), .B(G107), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NAND2_X1  g418(.A1(new_n580), .A2(new_n292), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n350), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n350), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT94), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n608), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n354), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n611), .A2(new_n614), .A3(new_n349), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n360), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n358), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n605), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n410), .A2(KEYINPUT92), .A3(new_n415), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT92), .B1(new_n410), .B2(new_n415), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI211_X1 g437(.A(G902), .B(new_n572), .C1(new_n567), .C2(new_n570), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n531), .B1(new_n624), .B2(new_n560), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n592), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n620), .A2(new_n623), .A3(new_n626), .A4(new_n457), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  NOR2_X1   g443(.A1(new_n334), .A2(G900), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(G902), .A3(new_n450), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n633), .A2(new_n634), .A3(new_n452), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(KEYINPUT97), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n601), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n619), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(new_n626), .A3(new_n296), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT98), .B(G128), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G30));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n638), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT39), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT40), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n290), .A2(new_n266), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n254), .A2(new_n255), .A3(new_n263), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(G902), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n294), .B(new_n295), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n526), .A2(new_n527), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n648), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n418), .A2(new_n419), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n528), .A3(new_n449), .A4(new_n619), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n204), .ZN(G45));
  NAND3_X1  g475(.A1(new_n626), .A2(new_n296), .A3(new_n640), .ZN(new_n662));
  INV_X1    g476(.A(new_n586), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n644), .C1(new_n621), .C2(new_n622), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n202), .ZN(G48));
  NAND2_X1  g480(.A1(new_n587), .A2(new_n593), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n562), .A2(KEYINPUT81), .B1(new_n554), .B2(new_n555), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(new_n566), .B1(new_n569), .B2(new_n543), .ZN(new_n669));
  OAI21_X1  g483(.A(G469), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n531), .A3(new_n574), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n574), .A3(KEYINPUT100), .A4(new_n531), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n296), .A2(new_n673), .A3(new_n362), .A4(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT41), .B(G113), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NAND3_X1  g492(.A1(new_n593), .A2(new_n600), .A3(new_n599), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n675), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n197), .ZN(G18));
  NAND3_X1  g495(.A1(new_n673), .A2(new_n530), .A3(new_n674), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n296), .A2(new_n640), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n458), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n195), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n530), .A2(new_n449), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n686), .B1(new_n623), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n592), .A2(new_n598), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n658), .A2(new_n689), .A3(KEYINPUT103), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n580), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n257), .B1(new_n256), .B2(new_n269), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n249), .A2(KEYINPUT70), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT101), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n253), .A2(new_n258), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n266), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n290), .A2(new_n263), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT102), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n698), .A2(new_n703), .A3(new_n700), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n287), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n692), .B1(new_n705), .B2(new_n283), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n673), .A2(new_n674), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n707), .A2(new_n456), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n691), .A2(new_n362), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  INV_X1    g524(.A(new_n664), .ZN(new_n711));
  INV_X1    g525(.A(new_n682), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n706), .A2(new_n711), .A3(new_n712), .A4(new_n640), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  NOR3_X1   g528(.A1(new_n533), .A2(KEYINPUT104), .A3(G902), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n549), .B(new_n715), .C1(new_n558), .C2(new_n544), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(new_n560), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n532), .B1(new_n718), .B2(new_n574), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n529), .B1(new_n590), .B2(new_n591), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT32), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n292), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n280), .A2(new_n725), .A3(new_n295), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n362), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n727), .B1(new_n726), .B2(new_n362), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n723), .B(new_n711), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n296), .A2(new_n719), .A3(new_n362), .A4(new_n720), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n722), .B1(new_n732), .B2(new_n664), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT106), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n732), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n639), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n621), .A2(new_n622), .A3(new_n586), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(KEYINPUT107), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n744), .B(KEYINPUT43), .C1(new_n658), .C2(new_n586), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n619), .B1(new_n292), .B2(new_n580), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n743), .A2(new_n745), .A3(KEYINPUT44), .A4(new_n746), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n533), .A2(new_n187), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n533), .B1(new_n559), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n549), .B(KEYINPUT45), .C1(new_n558), .C2(new_n544), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n574), .B1(new_n755), .B2(KEYINPUT46), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n757), .B(new_n751), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n531), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n646), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n720), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  AOI21_X1  g578(.A(new_n263), .B1(new_n256), .B2(new_n269), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n276), .A2(new_n266), .A3(new_n254), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(new_n286), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n282), .B1(new_n767), .B2(new_n700), .ZN(new_n768));
  AOI22_X1  g582(.A1(KEYINPUT32), .A2(new_n768), .B1(new_n279), .B2(G472), .ZN(new_n769));
  INV_X1    g583(.A(new_n362), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n294), .A3(new_n770), .A4(new_n720), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n664), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n759), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n531), .B(new_n773), .C1(new_n756), .C2(new_n758), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  AND2_X1   g592(.A1(new_n743), .A2(new_n745), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n706), .A2(new_n362), .A3(new_n452), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n656), .A2(new_n528), .A3(new_n707), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n775), .A2(new_n776), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n670), .A2(new_n574), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n531), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n720), .A3(new_n779), .A4(new_n780), .ZN(new_n788));
  NOR2_X1   g602(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n673), .A2(new_n674), .A3(new_n720), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT114), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n673), .A2(new_n793), .A3(new_n674), .A4(new_n720), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n452), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n653), .A2(new_n770), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n623), .A3(new_n586), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n784), .A2(new_n788), .A3(new_n790), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n704), .A2(new_n287), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n703), .B1(new_n698), .B2(new_n700), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n283), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n580), .A3(new_n640), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n779), .A2(new_n796), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n743), .A2(new_n745), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT115), .B1(new_n806), .B2(new_n795), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n799), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n811), .B2(KEYINPUT51), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n796), .A2(new_n587), .A3(new_n797), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(G952), .A3(new_n334), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n779), .A2(new_n780), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n712), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n805), .A2(new_n807), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n726), .A2(new_n362), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n728), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n817), .B2(new_n820), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n811), .B2(KEYINPUT51), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n826), .B(new_n827), .C1(new_n830), .C2(new_n799), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n812), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n581), .A2(new_n587), .A3(new_n593), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n577), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n623), .A2(new_n626), .A3(new_n457), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n594), .B(KEYINPUT109), .C1(new_n363), .C2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n709), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n675), .B1(new_n667), .B2(new_n679), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n684), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n623), .A2(new_n449), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n627), .B1(new_n597), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n619), .A2(new_n653), .A3(new_n644), .A4(new_n719), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n658), .A2(new_n689), .A3(KEYINPUT103), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT103), .B1(new_n658), .B2(new_n689), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n683), .A2(new_n576), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n639), .B2(new_n711), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n713), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n849), .A2(new_n713), .A3(new_n851), .A4(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n447), .A2(new_n448), .A3(new_n644), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(G475), .B2(new_n414), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n600), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n720), .A2(new_n859), .A3(new_n575), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT110), .B1(new_n683), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n528), .B1(new_n526), .B2(new_n527), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n600), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n862), .A2(new_n625), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n296), .A4(new_n640), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n739), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n803), .A2(new_n664), .A3(new_n721), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT111), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n861), .A2(new_n866), .B1(new_n738), .B2(new_n639), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  INV_X1    g686(.A(new_n721), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n706), .A2(new_n711), .A3(new_n640), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n845), .A2(new_n856), .A3(new_n876), .A4(new_n736), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT53), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n872), .A2(new_n874), .A3(new_n867), .A4(new_n739), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n872), .B1(new_n871), .B2(new_n874), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n842), .A2(new_n839), .A3(new_n684), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n709), .A3(new_n837), .A4(new_n835), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n736), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n854), .A2(KEYINPUT112), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n878), .B(KEYINPUT54), .C1(new_n886), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n885), .B1(new_n731), .B2(new_n733), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n884), .A2(new_n887), .A3(new_n888), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n877), .A2(new_n885), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n890), .B1(KEYINPUT54), .B2(new_n894), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n832), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n586), .A2(new_n532), .A3(new_n529), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(KEYINPUT49), .B2(new_n786), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(KEYINPUT49), .B2(new_n786), .ZN(new_n899));
  INV_X1    g713(.A(new_n656), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n623), .A4(new_n797), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(G75));
  NAND3_X1  g716(.A1(new_n894), .A2(G902), .A3(new_n505), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n495), .B(KEYINPUT119), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n502), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n334), .A2(G952), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n751), .B(KEYINPUT57), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT54), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n892), .A2(new_n893), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n892), .B2(new_n893), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n571), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n894), .A2(G902), .A3(new_n754), .A4(new_n753), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n894), .A2(G902), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n397), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n910), .ZN(G60));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n584), .B1(new_n895), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n584), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n914), .B2(new_n915), .ZN(new_n932));
  INV_X1    g746(.A(new_n910), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n930), .A2(new_n934), .ZN(G63));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n297), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n892), .B2(new_n893), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n616), .A2(new_n617), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n359), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n933), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n936), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n892), .A2(new_n893), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n359), .B1(new_n945), .B2(new_n937), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n933), .A4(new_n940), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(G66));
  OAI21_X1  g762(.A(G953), .B1(new_n455), .B2(new_n500), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n845), .B2(G953), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n905), .B1(G898), .B2(new_n334), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n284), .B(KEYINPUT122), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(new_n393), .Z(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n955), .B(new_n956), .Z(new_n957));
  INV_X1    g771(.A(new_n363), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n862), .A2(new_n625), .A3(new_n646), .ZN(new_n959));
  INV_X1    g773(.A(new_n841), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n958), .B(new_n959), .C1(new_n960), .C2(new_n587), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n777), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n761), .B1(new_n747), .B2(new_n748), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n750), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n803), .A2(new_n664), .A3(new_n682), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n641), .B1(new_n662), .B2(new_n664), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n713), .A2(new_n851), .A3(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n660), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n657), .A2(new_n659), .ZN(new_n973));
  INV_X1    g787(.A(new_n969), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT123), .B1(new_n713), .B2(new_n851), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n973), .B(new_n971), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n970), .A2(new_n978), .A3(new_n971), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n972), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n953), .B(new_n957), .C1(new_n980), .C2(G953), .ZN(new_n981));
  INV_X1    g795(.A(G900), .ZN(new_n982));
  OAI21_X1  g796(.A(G953), .B1(new_n541), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n957), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n972), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n987), .B2(new_n334), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n968), .A2(new_n969), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n691), .A2(new_n820), .A3(new_n760), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n777), .A2(new_n739), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n736), .A2(new_n989), .A3(new_n763), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n630), .B1(new_n993), .B2(new_n334), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT125), .B1(new_n994), .B2(new_n957), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n981), .B(new_n983), .C1(new_n988), .C2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n957), .B1(new_n980), .B2(G953), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n731), .A2(new_n733), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT106), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n733), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n992), .A2(new_n763), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n989), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n334), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n630), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n953), .B1(new_n1007), .B2(new_n984), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n998), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n983), .B1(new_n1009), .B2(new_n981), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n997), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT63), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT126), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n993), .B2(new_n883), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n266), .B(new_n290), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n987), .B2(new_n883), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n649), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1013), .B1(new_n699), .B2(new_n277), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n878), .B(new_n1021), .C1(new_n886), .C2(new_n889), .ZN(new_n1022));
  AND4_X1   g836(.A1(new_n933), .A2(new_n1018), .A3(new_n1020), .A4(new_n1022), .ZN(G57));
endmodule


