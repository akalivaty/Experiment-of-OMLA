

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n369), .B(n313), .ZN(n314) );
  XOR2_X1 U326 ( .A(G162GAT), .B(G218GAT), .Z(n359) );
  XNOR2_X1 U327 ( .A(n319), .B(n318), .ZN(n326) );
  XNOR2_X1 U328 ( .A(n396), .B(n395), .ZN(n571) );
  XNOR2_X1 U329 ( .A(n394), .B(KEYINPUT98), .ZN(n395) );
  XNOR2_X1 U330 ( .A(n449), .B(KEYINPUT38), .ZN(n504) );
  AND2_X1 U331 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  NOR2_X1 U332 ( .A1(n536), .A2(n524), .ZN(n470) );
  XNOR2_X1 U333 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n459) );
  INV_X1 U334 ( .A(KEYINPUT31), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n365), .B(n293), .ZN(n366) );
  INV_X1 U336 ( .A(G85GAT), .ZN(n318) );
  XNOR2_X1 U337 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U338 ( .A(n367), .B(n366), .ZN(n368) );
  INV_X1 U339 ( .A(KEYINPUT119), .ZN(n474) );
  INV_X1 U340 ( .A(KEYINPUT26), .ZN(n394) );
  XNOR2_X1 U341 ( .A(n326), .B(n380), .ZN(n323) );
  XNOR2_X1 U342 ( .A(n372), .B(n408), .ZN(n373) );
  XNOR2_X1 U343 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  XNOR2_X1 U344 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U345 ( .A(n374), .B(n373), .ZN(n376) );
  XNOR2_X1 U346 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U347 ( .A(n325), .B(n324), .ZN(n453) );
  NOR2_X1 U348 ( .A1(n528), .A2(n477), .ZN(n568) );
  XOR2_X1 U349 ( .A(n453), .B(KEYINPUT41), .Z(n542) );
  INV_X1 U350 ( .A(KEYINPUT104), .ZN(n450) );
  XNOR2_X1 U351 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n478) );
  XNOR2_X1 U352 ( .A(n450), .B(G50GAT), .ZN(n451) );
  XNOR2_X1 U353 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U354 ( .A(n452), .B(n451), .ZN(G1331GAT) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n294) );
  XNOR2_X1 U356 ( .A(n294), .B(G29GAT), .ZN(n295) );
  XOR2_X1 U357 ( .A(n295), .B(KEYINPUT8), .Z(n297) );
  XNOR2_X1 U358 ( .A(G43GAT), .B(G50GAT), .ZN(n296) );
  XOR2_X1 U359 ( .A(n297), .B(n296), .Z(n327) );
  XOR2_X1 U360 ( .A(G15GAT), .B(G1GAT), .Z(n348) );
  XOR2_X1 U361 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n299) );
  NAND2_X1 U362 ( .A1(G229GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U363 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U364 ( .A(n348), .B(n300), .Z(n301) );
  XNOR2_X1 U365 ( .A(n327), .B(n301), .ZN(n305) );
  XOR2_X1 U366 ( .A(G113GAT), .B(G197GAT), .Z(n303) );
  XNOR2_X1 U367 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n302) );
  XNOR2_X1 U368 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U369 ( .A(n305), .B(n304), .Z(n307) );
  XOR2_X1 U370 ( .A(G22GAT), .B(G141GAT), .Z(n360) );
  XOR2_X1 U371 ( .A(G169GAT), .B(G8GAT), .Z(n400) );
  XNOR2_X1 U372 ( .A(n360), .B(n400), .ZN(n306) );
  XNOR2_X1 U373 ( .A(n307), .B(n306), .ZN(n573) );
  XNOR2_X1 U374 ( .A(KEYINPUT69), .B(n573), .ZN(n567) );
  INV_X1 U375 ( .A(n567), .ZN(n465) );
  XOR2_X1 U376 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n309) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .Z(n344) );
  XOR2_X1 U378 ( .A(G176GAT), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U379 ( .A(n344), .B(n399), .ZN(n308) );
  XNOR2_X1 U380 ( .A(n309), .B(n308), .ZN(n315) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(G78GAT), .ZN(n310) );
  XNOR2_X1 U382 ( .A(n310), .B(G204GAT), .ZN(n369) );
  NAND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XOR2_X1 U384 ( .A(n315), .B(n314), .Z(n325) );
  XOR2_X1 U385 ( .A(KEYINPUT71), .B(G92GAT), .Z(n317) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(G106GAT), .ZN(n316) );
  XNOR2_X1 U387 ( .A(n317), .B(n316), .ZN(n319) );
  XOR2_X1 U388 ( .A(G71GAT), .B(G120GAT), .Z(n380) );
  XOR2_X1 U389 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n321) );
  XNOR2_X1 U390 ( .A(KEYINPUT74), .B(KEYINPUT70), .ZN(n320) );
  XOR2_X1 U391 ( .A(n321), .B(n320), .Z(n322) );
  NOR2_X1 U392 ( .A1(n465), .A2(n453), .ZN(n491) );
  XOR2_X1 U393 ( .A(n327), .B(n326), .Z(n337) );
  XOR2_X1 U394 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n329) );
  XNOR2_X1 U395 ( .A(KEYINPUT75), .B(KEYINPUT11), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U397 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n331) );
  XOR2_X1 U398 ( .A(G190GAT), .B(G134GAT), .Z(n381) );
  XNOR2_X1 U399 ( .A(n381), .B(n359), .ZN(n330) );
  XNOR2_X1 U400 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U401 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U402 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U404 ( .A(n337), .B(n336), .Z(n564) );
  INV_X1 U405 ( .A(n564), .ZN(n458) );
  XOR2_X1 U406 ( .A(KEYINPUT77), .B(n458), .Z(n548) );
  XNOR2_X1 U407 ( .A(KEYINPUT36), .B(n548), .ZN(n585) );
  XOR2_X1 U408 ( .A(G211GAT), .B(KEYINPUT12), .Z(n339) );
  XNOR2_X1 U409 ( .A(G22GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U410 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U411 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n341) );
  XNOR2_X1 U412 ( .A(G71GAT), .B(KEYINPUT80), .ZN(n340) );
  XNOR2_X1 U413 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U414 ( .A(n343), .B(n342), .Z(n350) );
  XOR2_X1 U415 ( .A(G127GAT), .B(n344), .Z(n346) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U418 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U419 ( .A(n350), .B(n349), .ZN(n358) );
  XOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n352) );
  XNOR2_X1 U421 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n351) );
  XNOR2_X1 U422 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G78GAT), .Z(n354) );
  XNOR2_X1 U424 ( .A(G155GAT), .B(KEYINPUT82), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U426 ( .A(n356), .B(n355), .Z(n357) );
  XOR2_X1 U427 ( .A(n358), .B(n357), .Z(n560) );
  INV_X1 U428 ( .A(n560), .ZN(n582) );
  XOR2_X1 U429 ( .A(n359), .B(G106GAT), .Z(n362) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(n360), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U432 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n364) );
  XNOR2_X1 U433 ( .A(KEYINPUT85), .B(KEYINPUT23), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U435 ( .A(n368), .B(KEYINPUT87), .Z(n374) );
  XNOR2_X1 U436 ( .A(n369), .B(KEYINPUT88), .ZN(n372) );
  XOR2_X1 U437 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n371) );
  XNOR2_X1 U438 ( .A(G197GAT), .B(G211GAT), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n408) );
  XNOR2_X1 U440 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n375) );
  XOR2_X1 U441 ( .A(n375), .B(KEYINPUT2), .Z(n435) );
  XNOR2_X1 U442 ( .A(n376), .B(n435), .ZN(n473) );
  XOR2_X1 U443 ( .A(KEYINPUT18), .B(G183GAT), .Z(n378) );
  XNOR2_X1 U444 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U446 ( .A(KEYINPUT84), .B(n379), .Z(n412) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U448 ( .A(G113GAT), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U449 ( .A(n382), .B(KEYINPUT0), .ZN(n436) );
  XNOR2_X1 U450 ( .A(n383), .B(n436), .ZN(n387) );
  XOR2_X1 U451 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n385) );
  NAND2_X1 U452 ( .A1(G227GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U454 ( .A(n387), .B(n386), .Z(n392) );
  XOR2_X1 U455 ( .A(G176GAT), .B(G99GAT), .Z(n389) );
  XNOR2_X1 U456 ( .A(G43GAT), .B(G15GAT), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U458 ( .A(G169GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U460 ( .A(n412), .B(n393), .Z(n537) );
  INV_X1 U461 ( .A(n537), .ZN(n528) );
  NAND2_X1 U462 ( .A1(n473), .A2(n528), .ZN(n396) );
  XOR2_X1 U463 ( .A(KEYINPUT96), .B(G204GAT), .Z(n398) );
  XNOR2_X1 U464 ( .A(G36GAT), .B(G92GAT), .ZN(n397) );
  XNOR2_X1 U465 ( .A(n398), .B(n397), .ZN(n404) );
  XOR2_X1 U466 ( .A(n399), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U467 ( .A(n400), .B(G190GAT), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U469 ( .A(n404), .B(n403), .Z(n406) );
  NAND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U472 ( .A(n407), .B(KEYINPUT95), .Z(n410) );
  XNOR2_X1 U473 ( .A(n408), .B(KEYINPUT97), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U475 ( .A(n412), .B(n411), .Z(n513) );
  XNOR2_X1 U476 ( .A(KEYINPUT27), .B(n513), .ZN(n442) );
  NAND2_X1 U477 ( .A1(n571), .A2(n442), .ZN(n417) );
  XOR2_X1 U478 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n415) );
  INV_X1 U479 ( .A(n513), .ZN(n524) );
  NOR2_X1 U480 ( .A1(n528), .A2(n524), .ZN(n413) );
  NOR2_X1 U481 ( .A1(n473), .A2(n413), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  NAND2_X1 U483 ( .A1(n417), .A2(n416), .ZN(n441) );
  XOR2_X1 U484 ( .A(KEYINPUT89), .B(KEYINPUT6), .Z(n419) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U487 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n421) );
  XNOR2_X1 U488 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U490 ( .A(n423), .B(n422), .Z(n428) );
  XOR2_X1 U491 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n425) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U494 ( .A(KEYINPUT91), .B(n426), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U496 ( .A(G162GAT), .B(G85GAT), .Z(n430) );
  XNOR2_X1 U497 ( .A(G29GAT), .B(G134GAT), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U499 ( .A(G148GAT), .B(G57GAT), .Z(n432) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(G120GAT), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U502 ( .A(n434), .B(n433), .Z(n438) );
  XOR2_X1 U503 ( .A(n436), .B(n435), .Z(n437) );
  XNOR2_X1 U504 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n440), .B(n439), .ZN(n510) );
  INV_X1 U506 ( .A(n510), .ZN(n522) );
  NAND2_X1 U507 ( .A1(n441), .A2(n522), .ZN(n445) );
  XOR2_X1 U508 ( .A(KEYINPUT28), .B(n473), .Z(n531) );
  INV_X1 U509 ( .A(n531), .ZN(n540) );
  NAND2_X1 U510 ( .A1(n510), .A2(n442), .ZN(n535) );
  NOR2_X1 U511 ( .A1(n540), .A2(n535), .ZN(n443) );
  NAND2_X1 U512 ( .A1(n443), .A2(n528), .ZN(n444) );
  NAND2_X1 U513 ( .A1(n445), .A2(n444), .ZN(n446) );
  XOR2_X1 U514 ( .A(KEYINPUT100), .B(n446), .Z(n489) );
  NOR2_X1 U515 ( .A1(n582), .A2(n489), .ZN(n447) );
  NAND2_X1 U516 ( .A1(n585), .A2(n447), .ZN(n448) );
  XNOR2_X1 U517 ( .A(n448), .B(KEYINPUT37), .ZN(n521) );
  NAND2_X1 U518 ( .A1(n491), .A2(n521), .ZN(n449) );
  NOR2_X1 U519 ( .A1(n504), .A2(n531), .ZN(n452) );
  INV_X1 U520 ( .A(n542), .ZN(n556) );
  NOR2_X1 U521 ( .A1(n556), .A2(n573), .ZN(n454) );
  XNOR2_X1 U522 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  NOR2_X1 U523 ( .A1(n455), .A2(n582), .ZN(n456) );
  XNOR2_X1 U524 ( .A(n456), .B(KEYINPUT111), .ZN(n457) );
  NOR2_X1 U525 ( .A1(n458), .A2(n457), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n460), .B(n459), .ZN(n467) );
  XOR2_X1 U527 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n462) );
  NAND2_X1 U528 ( .A1(n582), .A2(n585), .ZN(n461) );
  XNOR2_X1 U529 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U530 ( .A1(n463), .A2(n453), .ZN(n464) );
  NAND2_X1 U531 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U532 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U533 ( .A(KEYINPUT48), .ZN(n468) );
  XNOR2_X1 U534 ( .A(n469), .B(n468), .ZN(n536) );
  XNOR2_X1 U535 ( .A(n470), .B(KEYINPUT54), .ZN(n471) );
  NAND2_X1 U536 ( .A1(n471), .A2(n522), .ZN(n472) );
  XNOR2_X1 U537 ( .A(n472), .B(KEYINPUT64), .ZN(n570) );
  NOR2_X1 U538 ( .A1(n570), .A2(n473), .ZN(n476) );
  NAND2_X1 U539 ( .A1(n568), .A2(n548), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n568), .A2(n582), .ZN(n482) );
  XOR2_X1 U541 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(G183GAT), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(G1350GAT) );
  NAND2_X1 U544 ( .A1(n568), .A2(n542), .ZN(n486) );
  XOR2_X1 U545 ( .A(G176GAT), .B(KEYINPUT56), .Z(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  NOR2_X1 U549 ( .A1(n548), .A2(n560), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U551 ( .A1(n489), .A2(n488), .ZN(n490) );
  XOR2_X1 U552 ( .A(KEYINPUT101), .B(n490), .Z(n508) );
  NAND2_X1 U553 ( .A1(n491), .A2(n508), .ZN(n499) );
  NOR2_X1 U554 ( .A1(n522), .A2(n499), .ZN(n492) );
  XOR2_X1 U555 ( .A(G1GAT), .B(n492), .Z(n493) );
  XNOR2_X1 U556 ( .A(KEYINPUT34), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U557 ( .A1(n524), .A2(n499), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(n494), .Z(n495) );
  XNOR2_X1 U559 ( .A(G8GAT), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U560 ( .A1(n528), .A2(n499), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U563 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NOR2_X1 U564 ( .A1(n531), .A2(n499), .ZN(n500) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U566 ( .A1(n504), .A2(n522), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n504), .A2(n524), .ZN(n503) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n503), .Z(G1329GAT) );
  NOR2_X1 U571 ( .A1(n504), .A2(n528), .ZN(n505) );
  XOR2_X1 U572 ( .A(KEYINPUT40), .B(n505), .Z(n506) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n512) );
  NAND2_X1 U575 ( .A1(n542), .A2(n573), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n507), .B(KEYINPUT105), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n520), .A2(n508), .ZN(n509) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n509), .Z(n517) );
  NAND2_X1 U579 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n513), .A2(n517), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n514), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(G71GAT), .B(KEYINPUT107), .Z(n516) );
  NAND2_X1 U584 ( .A1(n537), .A2(n517), .ZN(n515) );
  XNOR2_X1 U585 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U587 ( .A1(n540), .A2(n517), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n521), .A2(n520), .ZN(n530) );
  NOR2_X1 U590 ( .A1(n522), .A2(n530), .ZN(n523) );
  XOR2_X1 U591 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U592 ( .A1(n524), .A2(n530), .ZN(n526) );
  XNOR2_X1 U593 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U596 ( .A1(n528), .A2(n530), .ZN(n529) );
  XOR2_X1 U597 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U598 ( .A1(n531), .A2(n530), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n553) );
  NAND2_X1 U603 ( .A1(n537), .A2(n553), .ZN(n538) );
  XOR2_X1 U604 ( .A(KEYINPUT113), .B(n538), .Z(n539) );
  NOR2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n549), .A2(n567), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U609 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n546) );
  NAND2_X1 U612 ( .A1(n549), .A2(n582), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G127GAT), .B(n547), .Z(G1342GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U618 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U619 ( .A1(n571), .A2(n553), .ZN(n563) );
  NOR2_X1 U620 ( .A1(n573), .A2(n563), .ZN(n554) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n554), .Z(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT116), .B(n555), .ZN(G1344GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n563), .ZN(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n563), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT118), .B(n565), .Z(n566) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(n569), .ZN(G1348GAT) );
  INV_X1 U635 ( .A(n570), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n579) );
  NOR2_X1 U637 ( .A1(n573), .A2(n579), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U640 ( .A(n576), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U644 ( .A(n579), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n586), .A2(n453), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT125), .Z(n584) );
  NAND2_X1 U648 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

