//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n446, new_n450, new_n451, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n642, new_n644, new_n645, new_n646, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1269, new_n1270;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT68), .B(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n450));
  AND2_X1   g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  NAND2_X1  g027(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT71), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT72), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AND3_X1   g052(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G137), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(new_n462), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n472), .A2(new_n477), .A3(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n466), .A2(new_n467), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n485), .A2(KEYINPUT73), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(KEYINPUT73), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(G136), .A3(new_n462), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(G124), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n486), .A2(new_n487), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(new_n462), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n499), .B2(G124), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT74), .A3(new_n489), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(G162));
  INV_X1    g077(.A(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT3), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n465), .A2(G2104), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n504), .A2(new_n505), .A3(G138), .A4(new_n462), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT75), .B(G114), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n462), .ZN(new_n512));
  NAND2_X1  g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT4), .A2(G138), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(G2105), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n485), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G651), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT5), .B(G543), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n532), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT76), .B1(new_n525), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G88), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n532), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G303));
  INV_X1    g119(.A(G303), .ZN(G166));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT77), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT7), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n531), .A2(G51), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n535), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G168));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n535), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n536), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(new_n528), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n557), .A2(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n534), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n528), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n531), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n539), .A2(G81), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT78), .Z(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n522), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT79), .B(new_n573), .C1(new_n522), .C2(new_n574), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(G651), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n530), .ZN(new_n580));
  NOR2_X1   g155(.A1(KEYINPUT6), .A2(G651), .ZN(new_n581));
  OAI211_X1 g156(.A(G53), .B(G543), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n531), .A2(new_n584), .A3(G53), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n583), .A2(new_n585), .B1(new_n539), .B2(G91), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n579), .A2(new_n586), .ZN(G299));
  XNOR2_X1  g162(.A(G171), .B(KEYINPUT80), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  NAND2_X1  g164(.A1(new_n531), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n536), .ZN(G288));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n555), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n531), .A2(KEYINPUT83), .A3(G48), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n596), .A2(new_n597), .B1(G86), .B2(new_n539), .ZN(new_n598));
  OAI21_X1  g173(.A(G61), .B1(new_n520), .B2(new_n521), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(KEYINPUT81), .B1(G73), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n601), .B(G61), .C1(new_n520), .C2(new_n521), .ZN(new_n602));
  AOI211_X1 g177(.A(KEYINPUT82), .B(new_n528), .C1(new_n600), .C2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n604), .B1(new_n607), .B2(G651), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n603), .B2(new_n608), .ZN(G305));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  INV_X1    g185(.A(G47), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n536), .A2(new_n610), .B1(new_n555), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n528), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n612), .A2(new_n614), .ZN(G290));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n539), .A2(new_n616), .A3(G92), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT84), .B1(new_n536), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n534), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n528), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(G79), .A2(G543), .ZN(new_n626));
  INV_X1    g201(.A(G66), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n522), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT85), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n625), .A2(new_n629), .B1(G54), .B2(new_n531), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n622), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  XOR2_X1   g208(.A(G171), .B(KEYINPUT80), .Z(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(G868), .B2(new_n634), .ZN(G284));
  AOI21_X1  g210(.A(new_n633), .B1(G868), .B2(new_n634), .ZN(G321));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NAND2_X1  g212(.A1(G299), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(G168), .ZN(G297));
  OAI21_X1  g214(.A(new_n638), .B1(new_n637), .B2(G168), .ZN(G280));
  INV_X1    g215(.A(new_n632), .ZN(new_n641));
  INV_X1    g216(.A(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G860), .ZN(G148));
  OAI21_X1  g218(.A(KEYINPUT86), .B1(new_n566), .B2(G868), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n632), .A2(G559), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n645), .A2(new_n637), .ZN(new_n646));
  MUX2_X1   g221(.A(new_n644), .B(KEYINPUT86), .S(new_n646), .Z(G323));
  XNOR2_X1  g222(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g223(.A1(new_n498), .A2(G2105), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n499), .A2(G123), .ZN(new_n651));
  OR2_X1    g226(.A1(G99), .A2(G2105), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n652), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(G2096), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT87), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT12), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n657), .A3(new_n662), .ZN(G156));
  INV_X1    g238(.A(KEYINPUT14), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2427), .B(G2438), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2430), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT15), .B(G2435), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n667), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT16), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G14), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(G2072), .A2(G2078), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n444), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2067), .B(G2678), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n689), .A3(new_n685), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n683), .B(KEYINPUT17), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n690), .B(new_n681), .C1(new_n691), .C2(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n685), .A3(new_n680), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G2100), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT89), .B(G2096), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G227));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1956), .B(G2474), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1961), .B(G1966), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT20), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n700), .A2(new_n701), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n699), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n699), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(G1981), .B(G1986), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n710), .B(new_n714), .ZN(G229));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT91), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(KEYINPUT91), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G35), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n495), .A2(new_n496), .ZN(new_n724));
  AOI21_X1  g299(.A(KEYINPUT74), .B1(new_n500), .B2(new_n489), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n716), .B(new_n723), .C1(new_n726), .C2(new_n720), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n720), .B1(new_n497), .B2(new_n501), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT29), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(G2090), .A3(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n727), .A2(new_n729), .A3(KEYINPUT100), .A4(G2090), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1996), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n499), .B2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n649), .A2(G141), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n717), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n717), .A2(G32), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(KEYINPUT27), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n743), .A2(KEYINPUT27), .A3(new_n745), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n735), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n720), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(G116), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G2105), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n649), .B2(G140), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n499), .A2(KEYINPUT96), .A3(G128), .ZN(new_n756));
  AOI21_X1  g331(.A(KEYINPUT96), .B1(new_n499), .B2(G128), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n751), .B1(new_n758), .B2(G29), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G2067), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(G2067), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n743), .A2(KEYINPUT27), .A3(new_n745), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n763), .A2(new_n746), .A3(G1996), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n641), .A2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G4), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1348), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n765), .B(G1348), .C1(G4), .C2(G16), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT24), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G34), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n720), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G160), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n717), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2084), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n764), .A2(new_n768), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n762), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n717), .A2(G33), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n649), .A2(G139), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n781));
  NAND3_X1  g356(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OAI21_X1  g360(.A(G2105), .B1(new_n785), .B2(KEYINPUT98), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(KEYINPUT98), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n779), .B1(new_n788), .B2(new_n717), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2072), .ZN(new_n790));
  INV_X1    g365(.A(G299), .ZN(new_n791));
  INV_X1    g366(.A(G16), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G20), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT101), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n793), .A2(G1956), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(G1956), .B1(new_n793), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n792), .A2(G5), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G171), .B2(new_n792), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n797), .B(new_n798), .C1(new_n801), .C2(G1961), .ZN(new_n802));
  INV_X1    g377(.A(G28), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT30), .ZN(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n803), .B2(KEYINPUT30), .ZN(new_n805));
  OR2_X1    g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  NAND2_X1  g381(.A1(KEYINPUT31), .A2(G11), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(G16), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n565), .B2(new_n792), .ZN(new_n810));
  INV_X1    g385(.A(G1341), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n801), .A2(G1961), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n792), .A2(G21), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G168), .B2(new_n792), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n654), .A2(new_n721), .B1(G1966), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(G1966), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n721), .A2(G27), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G164), .B2(new_n721), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G2078), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n813), .A2(new_n814), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n790), .A2(new_n802), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n727), .A2(new_n729), .ZN(new_n825));
  INV_X1    g400(.A(G2090), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n734), .A2(new_n778), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n538), .A2(G16), .A3(new_n543), .ZN(new_n831));
  INV_X1    g406(.A(G1971), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n792), .A2(G22), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(G305), .A2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT32), .B(G1981), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT94), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n792), .A2(G6), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n792), .A2(G23), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G288), .B2(G16), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g420(.A(KEYINPUT33), .B(new_n842), .C1(G288), .C2(G16), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G1976), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  OAI21_X1  g425(.A(G1976), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n836), .A2(new_n841), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n837), .A2(new_n840), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n839), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n830), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n836), .A2(new_n852), .A3(new_n841), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n858), .A2(KEYINPUT95), .A3(new_n855), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n829), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n853), .A2(new_n830), .A3(new_n856), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT95), .B1(new_n858), .B2(new_n855), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT34), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n720), .A2(G25), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n649), .A2(G131), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n499), .A2(G119), .ZN(new_n866));
  OR2_X1    g441(.A1(G95), .A2(G2105), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n867), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n864), .B1(new_n869), .B2(new_n721), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G1991), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT92), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  MUX2_X1   g450(.A(G24), .B(G290), .S(G16), .Z(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT93), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(KEYINPUT93), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G1986), .ZN(new_n880));
  INV_X1    g455(.A(G1986), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n881), .A3(new_n878), .ZN(new_n882));
  AOI211_X1 g457(.A(new_n874), .B(new_n875), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n860), .A2(new_n863), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT36), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n860), .A2(new_n886), .A3(new_n863), .A4(new_n883), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n828), .B1(new_n885), .B2(new_n887), .ZN(G311));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n885), .A2(new_n887), .ZN(new_n890));
  INV_X1    g465(.A(new_n828), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(KEYINPUT102), .B(new_n828), .C1(new_n885), .C2(new_n887), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G150));
  INV_X1    g469(.A(G93), .ZN(new_n895));
  INV_X1    g470(.A(G55), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n536), .A2(new_n895), .B1(new_n555), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n534), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(new_n528), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n897), .B2(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G860), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT37), .Z(new_n906));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(new_n565), .A3(new_n903), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n565), .A2(new_n900), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT104), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT38), .Z(new_n915));
  NOR2_X1   g490(.A1(new_n632), .A2(new_n642), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n907), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G860), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n917), .A2(new_n918), .A3(new_n907), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n906), .B1(new_n921), .B2(new_n922), .ZN(G145));
  NAND2_X1  g498(.A1(new_n726), .A2(G160), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  NAND2_X1  g500(.A1(G162), .A2(new_n774), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n655), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n654), .A3(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n741), .A2(new_n742), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n788), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n787), .B2(new_n784), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n939));
  INV_X1    g514(.A(G118), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(G2105), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n499), .B2(G130), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n649), .A2(G142), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(new_n661), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n758), .A2(new_n517), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n758), .A2(new_n517), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n869), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n869), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n946), .A2(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n933), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n948), .A2(new_n955), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n932), .B(new_n930), .C1(new_n960), .C2(new_n957), .ZN(new_n961));
  INV_X1    g536(.A(G37), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g539(.A(new_n914), .B(new_n645), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n641), .B2(G299), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n641), .A2(G299), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n632), .A2(KEYINPUT106), .A3(new_n791), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT41), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT41), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n968), .A3(new_n972), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n965), .A2(new_n970), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(KEYINPUT107), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  INV_X1    g553(.A(G288), .ZN(new_n979));
  XNOR2_X1  g554(.A(G303), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(G305), .B(G290), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n975), .A2(new_n976), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  OAI21_X1  g562(.A(G868), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n904), .A2(new_n637), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(G295));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n989), .ZN(G331));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g571(.A1(G168), .A2(G171), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n634), .B2(G168), .ZN(new_n998));
  INV_X1    g573(.A(new_n913), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n997), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G301), .B2(G286), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n911), .A2(new_n1003), .A3(new_n913), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n970), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n971), .A2(new_n1001), .A3(new_n973), .A4(new_n1004), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n982), .ZN(new_n1009));
  INV_X1    g584(.A(new_n982), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  AND4_X1   g586(.A1(new_n996), .A2(new_n1009), .A3(new_n962), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G37), .B1(new_n1008), .B2(new_n982), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n996), .B1(new_n1013), .B2(new_n1011), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n994), .B(new_n995), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n962), .A3(new_n1011), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(new_n996), .A3(new_n1011), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n992), .A4(new_n993), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1015), .A2(new_n1019), .ZN(G397));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n517), .A2(new_n1022), .A3(KEYINPUT45), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n517), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n517), .B2(new_n1023), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n472), .A2(G40), .A3(new_n477), .A4(new_n483), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1971), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n517), .B2(new_n1023), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n517), .A2(new_n1034), .A3(new_n1023), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT113), .B(G2090), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1021), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(G114), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(KEYINPUT75), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(KEYINPUT75), .ZN(new_n1044));
  OAI21_X1  g619(.A(G2105), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1045), .A2(new_n510), .B1(new_n485), .B2(new_n515), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n1046), .B2(new_n508), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1025), .B(KEYINPUT111), .C1(new_n1047), .C2(new_n1028), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1031), .B1(new_n1048), .B2(new_n1024), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT116), .B(new_n1041), .C1(new_n1049), .C2(G1971), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1040), .A2(G8), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n538), .A2(G8), .A3(new_n543), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n538), .A2(KEYINPUT55), .A3(new_n543), .A4(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n517), .A2(new_n1023), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1031), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT114), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1062), .B(G8), .C1(new_n1031), .C2(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n598), .C1(new_n603), .C2(new_n608), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n596), .A2(new_n597), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n539), .A2(G86), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n528), .B1(new_n600), .B2(new_n602), .ZN(new_n1070));
  OAI21_X1  g645(.A(G1981), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(new_n1071), .A3(KEYINPUT49), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1064), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n979), .A2(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(G288), .B2(new_n848), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1078), .B(KEYINPUT115), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n482), .B1(new_n481), .B2(new_n462), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT72), .B(G2105), .C1(new_n480), .C2(new_n469), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(G40), .A3(new_n1047), .A4(new_n477), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1062), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1063), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1077), .B(new_n1079), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1076), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1064), .B2(new_n1077), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1037), .A2(KEYINPUT112), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n517), .A2(new_n1092), .A3(new_n1034), .A4(new_n1023), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1094), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1095));
  OAI211_X1 g670(.A(G8), .B(new_n1056), .C1(new_n1033), .C2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1058), .A2(new_n1090), .A3(KEYINPUT126), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1041), .B1(new_n1049), .B2(G1971), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1021), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1056), .B1(new_n1101), .B2(new_n1050), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT52), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(new_n1096), .A3(new_n1086), .A4(new_n1076), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1098), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1097), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G2078), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1049), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1094), .A2(new_n1036), .ZN(new_n1113));
  INV_X1    g688(.A(G1961), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT45), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1059), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n517), .A2(new_n1023), .A3(new_n1028), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1110), .A2(G2078), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1032), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1112), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1961), .B1(new_n1094), .B2(new_n1036), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1119), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1031), .A3(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1122), .A2(new_n1125), .A3(KEYINPUT123), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1111), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT124), .A3(new_n634), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n1049), .B2(new_n1108), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT123), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(G301), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(G40), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1082), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n476), .A2(KEYINPUT125), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n462), .B1(new_n476), .B2(KEYINPUT125), .ZN(new_n1138));
  AOI211_X1 g713(.A(new_n1135), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1030), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1111), .A2(new_n1140), .A3(new_n1115), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1141), .A2(new_n634), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1128), .A2(new_n1134), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1031), .A2(G2067), .A3(new_n1059), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1113), .B2(new_n767), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(new_n632), .ZN(new_n1149));
  AOI21_X1  g724(.A(G1348), .B1(new_n1094), .B2(new_n1036), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT118), .B(new_n641), .C1(new_n1150), .C2(new_n1147), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT56), .B(G2072), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1031), .B(new_n1153), .C1(new_n1048), .C2(new_n1024), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1956), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT57), .B1(G299), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n1158));
  AOI211_X1 g733(.A(KEYINPUT117), .B(new_n1158), .C1(new_n579), .C2(new_n586), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1154), .A2(new_n1155), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1149), .A2(new_n1151), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1030), .A2(new_n1032), .A3(new_n1152), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1035), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1032), .A2(new_n1163), .A3(new_n1037), .ZN(new_n1164));
  INV_X1    g739(.A(G1956), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1030), .A2(new_n735), .A3(new_n1032), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT58), .B(G1341), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n1083), .A2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n566), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n566), .B(new_n1177), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1150), .B2(new_n1147), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n632), .B1(new_n1148), .B2(KEYINPUT60), .ZN(new_n1184));
  NOR4_X1   g759(.A1(new_n1150), .A2(new_n641), .A3(new_n1182), .A4(new_n1147), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1167), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1187), .A2(new_n1188), .A3(KEYINPUT61), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n1160), .B2(new_n1168), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1186), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1169), .B1(new_n1181), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1133), .A2(G301), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1144), .B1(new_n1141), .B2(G171), .ZN(new_n1195));
  INV_X1    g770(.A(G2084), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1094), .A2(new_n1036), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(G1966), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1123), .B2(new_n1031), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(G8), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n1202));
  NOR2_X1   g777(.A1(G168), .A2(new_n1099), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1203), .A2(KEYINPUT51), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1099), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1203), .B(KEYINPUT121), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT51), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1204), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT122), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1205), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1212));
  AOI22_X1  g787(.A1(new_n1194), .A2(new_n1195), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1107), .A2(new_n1145), .A3(new_n1193), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1211), .A2(new_n1216), .A3(new_n1212), .ZN(new_n1217));
  AND2_X1   g792(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1219), .A2(KEYINPUT62), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1218), .A2(new_n1107), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1090), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1066), .ZN(new_n1223));
  NOR2_X1   g798(.A1(G288), .A2(G1976), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1076), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1064), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1222), .A2(new_n1096), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1201), .A2(G286), .ZN(new_n1228));
  NAND4_X1  g803(.A1(new_n1058), .A2(new_n1090), .A3(new_n1096), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT63), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g806(.A(G8), .B1(new_n1033), .B2(new_n1095), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1057), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1228), .A2(new_n1233), .A3(KEYINPUT63), .ZN(new_n1234));
  OR2_X1    g809(.A1(new_n1234), .A2(new_n1105), .ZN(new_n1235));
  AOI21_X1  g810(.A(new_n1227), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1214), .A2(new_n1221), .A3(new_n1236), .ZN(new_n1237));
  NOR3_X1   g812(.A1(new_n1031), .A2(new_n1047), .A3(new_n1028), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n758), .B(G2067), .ZN(new_n1239));
  INV_X1    g814(.A(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g815(.A(new_n934), .B(new_n735), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n869), .A2(new_n872), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n952), .A2(new_n873), .ZN(new_n1243));
  NAND4_X1  g818(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NOR2_X1   g819(.A1(G290), .A2(G1986), .ZN(new_n1245));
  NOR2_X1   g820(.A1(new_n1245), .A2(KEYINPUT110), .ZN(new_n1246));
  NAND2_X1  g821(.A1(G290), .A2(G1986), .ZN(new_n1247));
  XOR2_X1   g822(.A(new_n1246), .B(new_n1247), .Z(new_n1248));
  OAI21_X1  g823(.A(new_n1238), .B1(new_n1244), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1237), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1251));
  OAI22_X1  g826(.A1(new_n1251), .A2(new_n1243), .B1(G2067), .B2(new_n758), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1244), .A2(new_n1238), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1238), .A2(new_n1245), .ZN(new_n1254));
  XNOR2_X1  g829(.A(new_n1254), .B(KEYINPUT48), .ZN(new_n1255));
  AOI22_X1  g830(.A1(new_n1238), .A2(new_n1252), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1238), .B1(new_n1239), .B2(new_n934), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1238), .A2(new_n735), .ZN(new_n1258));
  XNOR2_X1  g833(.A(new_n1258), .B(KEYINPUT46), .ZN(new_n1259));
  NAND2_X1  g834(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g835(.A(new_n1260), .B(KEYINPUT47), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1256), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g839(.A1(new_n1256), .A2(new_n1261), .A3(KEYINPUT127), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1250), .A2(new_n1266), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g842(.A(G319), .B1(new_n677), .B2(new_n678), .ZN(new_n1269));
  NOR3_X1   g843(.A1(G229), .A2(G227), .A3(new_n1269), .ZN(new_n1270));
  OAI211_X1 g844(.A(new_n963), .B(new_n1270), .C1(new_n1014), .C2(new_n1012), .ZN(G225));
  INV_X1    g845(.A(G225), .ZN(G308));
endmodule


