//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT66), .Z(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n221), .B1(new_n206), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n223), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n202), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n227), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n219), .A2(new_n220), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G41), .A2(G45), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT67), .B1(new_n258), .B2(G1), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n260), .B(new_n261), .C1(G41), .C2(G45), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n257), .B1(new_n263), .B2(new_n209), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G77), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G222), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n271), .B1(new_n272), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n256), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n265), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n265), .A2(new_n278), .A3(KEYINPUT69), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G190), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n282), .A2(G200), .A3(new_n283), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n203), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(G150), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n267), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n288), .B1(new_n289), .B2(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n228), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n297), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n208), .B1(new_n261), .B2(G20), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(new_n208), .B2(new_n300), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n287), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n285), .A2(new_n286), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n285), .A2(new_n308), .A3(new_n311), .A4(new_n286), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n284), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n282), .A2(new_n316), .A3(new_n283), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n304), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n301), .ZN(new_n320));
  INV_X1    g0120(.A(new_n294), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n261), .A2(G20), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n320), .A2(new_n323), .B1(new_n299), .B2(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G58), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n210), .ZN(new_n327));
  OAI21_X1  g0127(.A(G20), .B1(new_n327), .B2(new_n202), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n290), .A2(G159), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT7), .B1(new_n333), .B2(new_n229), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n269), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT75), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n268), .A2(new_n229), .A3(new_n269), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n210), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT75), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT16), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n330), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n297), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n325), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT76), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n259), .A2(G232), .A3(new_n262), .A4(new_n256), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G223), .A2(G1698), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n209), .B2(G1698), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n270), .B1(G33), .B2(G87), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n257), .B(new_n351), .C1(new_n354), .C2(new_n256), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n254), .A2(new_n256), .A3(G274), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n209), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G223), .B2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n360), .B2(new_n333), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n357), .B1(new_n361), .B2(new_n277), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT77), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n363), .A3(new_n351), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n355), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n316), .B1(new_n314), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n346), .B1(new_n343), .B2(KEYINPUT75), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n338), .B(new_n210), .C1(new_n342), .C2(new_n335), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n297), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n343), .A2(new_n330), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n324), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n350), .A2(new_n367), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT18), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n355), .A2(G190), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n365), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n349), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n363), .B1(new_n362), .B2(new_n351), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n381), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n375), .A3(KEYINPUT17), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n350), .A2(new_n377), .A3(new_n392), .A4(new_n367), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n379), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n319), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT14), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n397));
  INV_X1    g0197(.A(G274), .ZN(new_n398));
  INV_X1    g0198(.A(new_n228), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n255), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(new_n254), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n209), .A2(new_n273), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n237), .A2(G1698), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n404), .C1(new_n331), .C2(new_n332), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n397), .A2(new_n402), .B1(new_n407), .B2(new_n277), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n263), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n259), .A2(KEYINPUT73), .A3(new_n262), .A4(new_n256), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G238), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n408), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n408), .B2(new_n412), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n396), .B(G169), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n410), .A2(G238), .A3(new_n411), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n401), .B1(new_n400), .B2(new_n254), .ZN(new_n418));
  AND4_X1   g0218(.A1(new_n401), .A2(new_n254), .A3(new_n256), .A4(G274), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G226), .A2(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n237), .B2(G1698), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n270), .B1(G33), .B2(G97), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n418), .A2(new_n419), .B1(new_n422), .B2(new_n256), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT13), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n408), .A2(new_n412), .A3(new_n413), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(G179), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n316), .B1(new_n424), .B2(new_n425), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n428), .A2(KEYINPUT74), .A3(new_n396), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT74), .ZN(new_n430));
  OAI21_X1  g0230(.A(G169), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(KEYINPUT14), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n427), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n300), .A2(new_n210), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT12), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n292), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n208), .B2(new_n291), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n301), .A2(G68), .A3(new_n322), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT11), .B1(new_n437), .B2(new_n297), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(G200), .B1(new_n414), .B2(new_n415), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n424), .A2(G190), .A3(new_n425), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n442), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT15), .B(G87), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n449));
  INV_X1    g0249(.A(G87), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT15), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT15), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G87), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n451), .A2(new_n453), .A3(KEYINPUT70), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n292), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n321), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n372), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n301), .A2(G77), .A3(new_n322), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G77), .B2(new_n299), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n211), .A2(G1698), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(G232), .B2(G1698), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n256), .B1(new_n463), .B2(new_n270), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G107), .B2(new_n270), .ZN(new_n465));
  INV_X1    g0265(.A(G244), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n257), .C1(new_n466), .C2(new_n263), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G200), .ZN(new_n468));
  INV_X1    g0268(.A(G190), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n461), .B(new_n468), .C1(new_n469), .C2(new_n467), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n461), .B1(new_n316), .B2(new_n467), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G179), .B2(new_n467), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n444), .A2(new_n447), .A3(new_n470), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n395), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G107), .ZN(new_n475));
  AND2_X1   g0275(.A1(KEYINPUT78), .A2(G97), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT78), .A2(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT6), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT6), .ZN(new_n479));
  AND2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  NOR2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n475), .B1(new_n342), .B2(new_n335), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI211_X1 g0287(.A(KEYINPUT79), .B(new_n475), .C1(new_n342), .C2(new_n335), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n297), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n299), .A2(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n261), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n299), .A2(new_n491), .A3(new_n228), .A4(new_n296), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n261), .A2(G45), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(KEYINPUT83), .B2(G41), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT83), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n252), .A3(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n506), .A2(new_n256), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G257), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n400), .A2(new_n501), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G244), .B(new_n273), .C1(new_n331), .C2(new_n332), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT80), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n270), .A2(new_n514), .A3(G244), .A4(new_n273), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT81), .A4(new_n516), .ZN(new_n520));
  OAI211_X1 g0320(.A(G250), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n512), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(KEYINPUT4), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT82), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n526), .A2(new_n527), .A3(new_n277), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(new_n526), .B2(new_n277), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n314), .B(new_n511), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n510), .B1(new_n526), .B2(new_n277), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n316), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n499), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n495), .B1(G190), .B2(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n526), .A2(new_n277), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT82), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n526), .A2(new_n527), .A3(new_n277), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n510), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n535), .B1(new_n539), .B2(new_n382), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n270), .A2(G244), .A3(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  OAI211_X1 g0342(.A(G238), .B(new_n273), .C1(new_n331), .C2(new_n332), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n277), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n501), .A2(new_n398), .ZN(new_n546));
  INV_X1    g0346(.A(G250), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n500), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n546), .A2(new_n256), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n451), .A2(new_n453), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT70), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n299), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n476), .A2(new_n477), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n293), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n229), .B1(new_n406), .B2(new_n558), .ZN(new_n561));
  OR2_X1    g0361(.A1(KEYINPUT78), .A2(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(KEYINPUT78), .A2(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n450), .A2(new_n475), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n270), .A2(new_n229), .A3(G68), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n568), .B2(new_n297), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n549), .B1(new_n544), .B2(new_n277), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G190), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n493), .A2(G87), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n552), .A2(new_n569), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n551), .A2(new_n316), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT85), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT85), .B1(new_n555), .B2(new_n556), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n493), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n570), .A2(new_n314), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT86), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n573), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n534), .A2(new_n540), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n270), .A2(new_n229), .A3(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n270), .A2(new_n589), .A3(new_n229), .A4(G87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n542), .A2(G20), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n229), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n475), .A2(KEYINPUT23), .A3(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n592), .B1(new_n591), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n297), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT25), .B1(new_n300), .B2(new_n475), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n475), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n604), .B1(G107), .B2(new_n493), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT88), .B(G294), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G33), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n606), .B(new_n608), .C1(new_n274), .C2(new_n547), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n277), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n507), .A2(G264), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n610), .A2(G190), .A3(new_n509), .A4(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n509), .A3(new_n611), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n601), .A2(new_n605), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n605), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n591), .A2(new_n597), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT24), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n598), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(new_n297), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n613), .A2(new_n316), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G179), .B2(new_n613), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n615), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n300), .A2(KEYINPUT87), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n299), .B2(G116), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n493), .A2(G116), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n229), .B(new_n522), .C1(new_n559), .C2(G33), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n296), .A2(new_n228), .B1(G20), .B2(new_n624), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT20), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(G33), .B1(new_n562), .B2(new_n563), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n522), .A2(new_n229), .ZN(new_n633));
  OAI211_X1 g0433(.A(KEYINPUT20), .B(new_n630), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n628), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n506), .A2(G270), .A3(new_n256), .ZN(new_n637));
  OAI211_X1 g0437(.A(G264), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n638));
  OAI211_X1 g0438(.A(G257), .B(new_n273), .C1(new_n331), .C2(new_n332), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n268), .A2(G303), .A3(new_n269), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n509), .B(new_n637), .C1(new_n641), .C2(new_n256), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(G200), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n469), .B2(new_n642), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n636), .A2(G169), .A3(new_n642), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n642), .A2(new_n314), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n645), .A2(new_n646), .B1(new_n647), .B2(new_n636), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n636), .A2(KEYINPUT21), .A3(G169), .A4(new_n642), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n644), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n474), .A2(new_n586), .A3(new_n651), .ZN(G372));
  INV_X1    g0452(.A(new_n318), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n349), .A2(new_n367), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(KEYINPUT18), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n392), .B1(new_n349), .B2(new_n367), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n447), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n444), .B1(new_n659), .B2(new_n472), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n391), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n661), .A2(new_n662), .B1(new_n310), .B2(new_n312), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n653), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n601), .A2(new_n605), .ZN(new_n666));
  INV_X1    g0466(.A(new_n613), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n314), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n621), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n648), .B2(new_n649), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n642), .A2(G169), .ZN(new_n672));
  INV_X1    g0472(.A(new_n627), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n299), .A2(new_n626), .A3(G116), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n673), .A2(new_n674), .B1(new_n624), .B2(new_n492), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n632), .A2(new_n633), .ZN(new_n677));
  INV_X1    g0477(.A(new_n630), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n679), .B2(new_n634), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n646), .B1(new_n672), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n647), .A2(new_n636), .ZN(new_n682));
  AND4_X1   g0482(.A1(new_n670), .A2(new_n681), .A3(new_n649), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n669), .B1(new_n671), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n581), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n615), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n534), .A3(new_n540), .A4(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n495), .A2(new_n573), .A3(new_n580), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n530), .A3(new_n689), .A4(new_n533), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(new_n580), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n573), .A2(new_n580), .A3(new_n583), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n583), .B1(new_n573), .B2(new_n580), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n534), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n687), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n474), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n665), .A2(new_n697), .ZN(G369));
  NOR2_X1   g0498(.A1(new_n671), .A2(new_n683), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n261), .A2(new_n229), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n680), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n699), .A2(KEYINPUT91), .A3(new_n707), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n650), .A2(new_n707), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n669), .B(new_n615), .C1(new_n620), .C2(new_n706), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n620), .A2(new_n622), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n716), .A2(KEYINPUT92), .A3(new_n705), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT92), .B1(new_n716), .B2(new_n705), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n648), .A2(new_n649), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n706), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n719), .A2(new_n725), .B1(new_n716), .B2(new_n706), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(G399));
  INV_X1    g0527(.A(new_n225), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n564), .A2(G116), .A3(new_n565), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n729), .A2(new_n731), .A3(new_n261), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n233), .B2(new_n729), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n733), .B(KEYINPUT28), .Z(new_n734));
  AND2_X1   g0534(.A1(new_n530), .A2(new_n533), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n585), .A3(new_n689), .A4(new_n499), .ZN(new_n736));
  INV_X1    g0536(.A(new_n580), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n688), .A2(new_n530), .A3(new_n533), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(KEYINPUT26), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n686), .B1(new_n716), .B2(new_n723), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n534), .A2(new_n540), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n736), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n706), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT94), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n696), .A2(new_n706), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n744), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n623), .A2(new_n650), .A3(new_n705), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(new_n585), .A3(new_n534), .A4(new_n540), .ZN(new_n752));
  AND4_X1   g0552(.A1(new_n570), .A2(new_n647), .A3(new_n611), .A4(new_n610), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n531), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(KEYINPUT30), .A3(new_n531), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n551), .A2(new_n314), .A3(new_n642), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n511), .B1(new_n528), .B2(new_n529), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n613), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n759), .B1(new_n761), .B2(KEYINPUT93), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n760), .A2(new_n763), .A3(new_n613), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n758), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n706), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n752), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(KEYINPUT93), .B1(new_n539), .B2(new_n667), .ZN(new_n770));
  INV_X1    g0570(.A(new_n759), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n764), .A3(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n756), .A2(new_n757), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(KEYINPUT31), .B1(new_n774), .B2(new_n705), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G330), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n750), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n734), .B1(new_n781), .B2(G1), .ZN(G364));
  AOI21_X1  g0582(.A(new_n228), .B1(G20), .B2(new_n316), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(G20), .A2(G179), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(new_n469), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G311), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n333), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n229), .A2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(new_n469), .A3(new_n382), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n789), .B(new_n793), .C1(G329), .C2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(new_n469), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G283), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n469), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n229), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n785), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n469), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n803), .A2(new_n607), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G303), .A2(new_n810), .B1(new_n812), .B2(G326), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n797), .A2(new_n800), .A3(new_n808), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n798), .A2(new_n475), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n809), .A2(new_n450), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G68), .C2(new_n806), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n270), .B1(new_n787), .B2(new_n326), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G77), .B2(new_n790), .ZN(new_n819));
  INV_X1    g0619(.A(G159), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n795), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n803), .A2(G97), .B1(new_n812), .B2(G50), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n817), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n784), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n223), .A2(G20), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n261), .B1(new_n826), .B2(G45), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n729), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(G13), .A2(G33), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(G20), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n783), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n233), .A2(new_n253), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n728), .A2(new_n270), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(new_n247), .C2(new_n253), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n728), .A2(new_n333), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G355), .B1(new_n624), .B2(new_n728), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n825), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n833), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n713), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n714), .A2(new_n830), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n713), .A2(G330), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT95), .ZN(G396));
  OR2_X1    g0648(.A1(new_n472), .A2(new_n705), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n470), .B1(new_n461), .B2(new_n706), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n472), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n746), .B(new_n852), .Z(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(new_n779), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n829), .B1(new_n853), .B2(new_n779), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n783), .A2(new_n831), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT96), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n829), .B1(new_n858), .B2(G77), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n832), .ZN(new_n860));
  INV_X1    g0660(.A(G283), .ZN(new_n861));
  INV_X1    g0661(.A(G303), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n805), .A2(new_n861), .B1(new_n811), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G87), .B2(new_n799), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n270), .B1(new_n796), .B2(G311), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G116), .A2(new_n790), .B1(new_n786), .B2(G294), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n803), .A2(G97), .B1(new_n810), .B2(G107), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(G143), .A2(new_n786), .B1(new_n790), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G137), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n870), .B2(new_n811), .C1(new_n289), .C2(new_n805), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT97), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT34), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n798), .A2(new_n210), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n333), .B(new_n874), .C1(G132), .C2(new_n796), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n803), .A2(G58), .B1(new_n810), .B2(G50), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n872), .A2(KEYINPUT34), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n868), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n859), .B(new_n860), .C1(new_n783), .C2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n856), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(G384));
  OR2_X1    g0682(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(G116), .A3(new_n230), .A4(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  NOR3_X1   g0686(.A1(new_n232), .A2(new_n272), .A3(new_n327), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT98), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(KEYINPUT98), .B1(G68), .B2(new_n201), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n261), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n368), .B1(new_n343), .B2(new_n330), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n324), .B1(new_n374), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n703), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n394), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n703), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n350), .A2(new_n377), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n389), .A2(new_n375), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n378), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n316), .B1(new_n385), .B2(new_n386), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n366), .A2(new_n314), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n894), .B1(new_n904), .B2(new_n703), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n349), .A2(new_n383), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n898), .B1(new_n657), .B2(new_n391), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n904), .A2(new_n375), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT100), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT100), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n654), .A2(new_n900), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n898), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n910), .B1(new_n916), .B2(new_n901), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n909), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n444), .A2(new_n705), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  INV_X1    g0724(.A(new_n895), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n384), .A2(new_n390), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(KEYINPUT18), .B2(new_n378), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n927), .B2(new_n393), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n901), .A2(new_n907), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n909), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n923), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n443), .B(new_n705), .C1(new_n433), .C2(new_n659), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n443), .A2(new_n705), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n416), .A2(new_n426), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT74), .B1(new_n428), .B2(new_n396), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n431), .A2(new_n430), .A3(KEYINPUT14), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n447), .B(new_n934), .C1(new_n938), .C2(new_n442), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n696), .A2(new_n706), .A3(new_n852), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n942), .B2(new_n849), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n930), .A2(new_n909), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n658), .A2(new_n703), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n932), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n745), .A2(new_n474), .A3(new_n748), .A4(new_n749), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n665), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n947), .B(new_n949), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n940), .A2(new_n852), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n766), .B1(new_n765), .B2(new_n706), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n774), .A2(new_n767), .B1(new_n586), .B2(new_n751), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n920), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT40), .B1(new_n930), .B2(new_n909), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(KEYINPUT40), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n776), .A2(new_n395), .A3(new_n473), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n777), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n959), .B2(new_n958), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n261), .B2(new_n826), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n950), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n892), .B1(new_n963), .B2(new_n964), .ZN(G367));
  XOR2_X1   g0765(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n809), .B2(new_n624), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT106), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n809), .A2(new_n624), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n969), .A2(KEYINPUT46), .B1(new_n806), .B2(new_n607), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n972));
  INV_X1    g0772(.A(G317), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n333), .B1(new_n795), .B2(new_n973), .C1(new_n559), .C2(new_n798), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G283), .A2(new_n790), .B1(new_n786), .B2(G303), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n475), .B2(new_n802), .C1(new_n792), .C2(new_n811), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n972), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n809), .A2(new_n326), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n802), .A2(new_n210), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(G159), .C2(new_n806), .ZN(new_n984));
  INV_X1    g0784(.A(new_n201), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n333), .B1(new_n985), .B2(new_n790), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n796), .A2(G137), .B1(new_n786), .B2(G150), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G77), .A2(new_n799), .B1(new_n812), .B2(G143), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n981), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT47), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n783), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n569), .A2(new_n572), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n705), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n580), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT101), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n685), .A2(new_n994), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(KEYINPUT101), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n833), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n835), .B1(new_n455), .B2(new_n728), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n837), .A2(new_n243), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n830), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n992), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n495), .A2(new_n705), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n534), .A2(new_n540), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n735), .A2(new_n495), .A3(new_n705), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n726), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n726), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1012), .A2(new_n1013), .B1(new_n721), .B2(KEYINPUT104), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n726), .A2(new_n1009), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(KEYINPUT102), .A3(KEYINPUT44), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT102), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT44), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n726), .A2(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT104), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n722), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1014), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1023), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT103), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n719), .B2(new_n725), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n714), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n713), .A3(G330), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n720), .A2(new_n724), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1031), .A2(new_n1034), .A3(new_n1032), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n779), .A3(new_n750), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n781), .B1(new_n1027), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n729), .B(KEYINPUT41), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n828), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1034), .A2(new_n1009), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT42), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n669), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n534), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n706), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT42), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1034), .A2(new_n1049), .A3(new_n1009), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1051), .A2(KEYINPUT43), .A3(new_n999), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT43), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1000), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n721), .A2(new_n1009), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1052), .A2(new_n721), .A3(new_n1009), .A4(new_n1056), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1005), .B1(new_n1043), .B2(new_n1061), .ZN(G387));
  NAND2_X1  g0862(.A1(new_n1038), .A2(new_n828), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G303), .A2(new_n790), .B1(new_n786), .B2(G317), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n792), .B2(new_n805), .C1(new_n788), .C2(new_n811), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n803), .A2(G283), .B1(new_n810), .B2(new_n607), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT112), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n798), .A2(new_n624), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n270), .B(new_n1074), .C1(G326), .C2(new_n796), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n575), .A2(new_n576), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n802), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n809), .A2(new_n272), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G150), .B2(new_n796), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT111), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n270), .B1(new_n791), .B2(new_n210), .C1(new_n208), .C2(new_n787), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G159), .A2(new_n812), .B1(new_n806), .B2(new_n321), .ZN(new_n1083));
  INV_X1    g0883(.A(G97), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n798), .ZN(new_n1085));
  OR4_X1    g0885(.A1(new_n1078), .A2(new_n1081), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n784), .B1(new_n1076), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n839), .A2(new_n731), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(G107), .B2(new_n225), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n240), .A2(G45), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT109), .Z(new_n1091));
  INV_X1    g0891(.A(new_n837), .ZN(new_n1092));
  AOI211_X1 g0892(.A(G45), .B(new_n731), .C1(G68), .C2(G77), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n294), .A2(G50), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1092), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1089), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n829), .B1(new_n1098), .B2(new_n835), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1087), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT113), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n719), .B2(new_n843), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1039), .A2(new_n729), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n781), .A2(new_n1038), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1063), .B1(new_n1102), .B2(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(G393));
  INV_X1    g0907(.A(new_n729), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1026), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1024), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1039), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1027), .A2(new_n1039), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n828), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n787), .A2(new_n820), .B1(new_n811), .B2(new_n289), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n333), .B1(new_n796), .B2(G143), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n294), .B2(new_n791), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n798), .A2(new_n450), .B1(new_n805), .B2(new_n201), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n802), .A2(new_n272), .B1(new_n809), .B2(new_n210), .ZN(new_n1122));
  OR4_X1    g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n787), .A2(new_n792), .B1(new_n811), .B2(new_n973), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT52), .ZN(new_n1125));
  INV_X1    g0925(.A(G294), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n333), .B1(new_n791), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G322), .B2(new_n796), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n815), .B1(G116), .B2(new_n803), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G283), .A2(new_n810), .B1(new_n806), .B2(G303), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n784), .B1(new_n1123), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1092), .A2(new_n250), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n835), .B1(new_n728), .B2(new_n564), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n830), .B(new_n1132), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1009), .B2(new_n843), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1114), .A2(new_n1115), .A3(new_n1136), .ZN(G390));
  AND3_X1   g0937(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n909), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n899), .B1(new_n349), .B2(new_n383), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n371), .A2(new_n374), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n376), .B1(new_n1140), .B2(new_n325), .ZN(new_n1141));
  AOI211_X1 g0941(.A(KEYINPUT76), .B(new_n324), .C1(new_n371), .C2(new_n374), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1143), .B2(new_n367), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n915), .A2(KEYINPUT37), .B1(new_n898), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n918), .B1(new_n1145), .B2(new_n910), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT39), .B1(new_n1146), .B2(new_n909), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n1138), .A2(new_n1147), .B1(new_n943), .B2(new_n923), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n923), .B1(new_n1146), .B2(new_n909), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n742), .A2(new_n706), .A3(new_n851), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n849), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1149), .B1(new_n1152), .B2(new_n941), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n953), .A2(new_n952), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1154), .A2(G330), .A3(new_n852), .A4(new_n940), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1148), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1156), .A2(new_n1157), .A3(new_n827), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n831), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1161), .A2(new_n790), .B1(G132), .B2(new_n786), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n795), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n803), .A2(G159), .B1(new_n812), .B2(G128), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n870), .B2(new_n805), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT53), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n809), .B2(new_n289), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n810), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1164), .B(new_n1166), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n270), .B1(new_n798), .B2(new_n201), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT116), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n802), .A2(new_n272), .B1(new_n787), .B2(new_n624), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT117), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n333), .B1(new_n795), .B2(new_n1126), .C1(new_n791), .C2(new_n559), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n805), .A2(new_n475), .B1(new_n811), .B2(new_n861), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n816), .A4(new_n874), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1170), .A2(new_n1172), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n829), .B1(new_n321), .B2(new_n858), .C1(new_n1178), .C2(new_n784), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT118), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n1159), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(KEYINPUT119), .B1(new_n1158), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1155), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1148), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1184), .B(new_n1181), .C1(new_n1189), .C2(new_n827), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n778), .A2(new_n474), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n948), .A2(new_n665), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n852), .C1(new_n769), .C2(new_n775), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n941), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1155), .A3(new_n1152), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT115), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1155), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n942), .A2(new_n849), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1195), .A2(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1194), .A2(new_n1155), .A3(KEYINPUT115), .A4(new_n1152), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1192), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n729), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1200), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1192), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(new_n1189), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1183), .B(new_n1190), .C1(new_n1203), .C2(new_n1209), .ZN(G378));
  NAND3_X1  g1010(.A1(new_n319), .A2(new_n304), .A3(new_n897), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n304), .A2(new_n897), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n313), .A2(new_n318), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n957), .B2(new_n777), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n956), .A2(new_n954), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT40), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n954), .B2(new_n920), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G330), .B(new_n1219), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1221), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n947), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1221), .A2(new_n947), .A3(new_n1226), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1220), .A2(new_n831), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n829), .B1(new_n858), .B2(new_n985), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G58), .A2(new_n799), .B1(new_n812), .B2(G116), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1084), .B2(new_n805), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n270), .A2(G41), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n861), .B2(new_n795), .C1(new_n475), .C2(new_n787), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1235), .A2(new_n1237), .A3(new_n983), .A4(new_n1079), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1077), .B2(new_n791), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT120), .Z(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT58), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT58), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G33), .A2(G41), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1236), .A2(G50), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G132), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n805), .A2(new_n1245), .B1(new_n811), .B2(new_n1163), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G150), .B2(new_n803), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G128), .A2(new_n786), .B1(new_n790), .B2(G137), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n809), .C2(new_n1160), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1250));
  INV_X1    g1050(.A(G124), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1243), .B1(new_n795), .B2(new_n1251), .C1(new_n820), .C2(new_n798), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1249), .B2(KEYINPUT59), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1244), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1241), .A2(new_n1242), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1233), .B1(new_n1255), .B2(new_n783), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1231), .A2(new_n828), .B1(new_n1232), .B2(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1221), .A2(new_n947), .A3(new_n1226), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n947), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1192), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n729), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1204), .A2(new_n1200), .A3(new_n1205), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1207), .B1(new_n1189), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1257), .B1(new_n1262), .B2(new_n1265), .ZN(G375));
  NAND4_X1  g1066(.A1(new_n1192), .A2(new_n1204), .A3(new_n1200), .A4(new_n1205), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1041), .B(KEYINPUT121), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1208), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n941), .A2(new_n831), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n829), .B1(new_n858), .B2(G68), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n809), .A2(new_n820), .B1(new_n811), .B2(new_n1245), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G50), .B2(new_n803), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n333), .B1(G137), .B2(new_n786), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n796), .A2(G128), .B1(G150), .B2(new_n790), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G58), .A2(new_n799), .B1(new_n806), .B2(new_n1161), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(G77), .A2(new_n799), .B1(new_n812), .B2(G294), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(G97), .A2(new_n810), .B1(new_n806), .B2(G116), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n270), .B1(G283), .B2(new_n786), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n796), .A2(G303), .B1(G107), .B2(new_n790), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1277), .B1(new_n1078), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1271), .B1(new_n1283), .B2(new_n783), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1206), .A2(new_n828), .B1(new_n1270), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1269), .A2(new_n1285), .ZN(G381));
  OR4_X1    g1086(.A1(G396), .A2(G381), .A3(G393), .A4(G384), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1136), .B1(new_n1027), .B2(new_n827), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1289), .B(new_n1005), .C1(new_n1043), .C2(new_n1061), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1181), .B1(new_n1189), .B2(new_n827), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1108), .B1(new_n1208), .B2(new_n1189), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  OR4_X1    g1095(.A1(G375), .A2(new_n1287), .A3(new_n1290), .A4(new_n1295), .ZN(G407));
  NAND2_X1  g1096(.A1(new_n704), .A2(G213), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G407), .B(G213), .C1(G375), .C2(new_n1299), .ZN(G409));
  AOI21_X1  g1100(.A(new_n1039), .B1(new_n1109), .B2(new_n1024), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1042), .B1(new_n1301), .B2(new_n780), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1061), .B1(new_n1302), .B2(new_n827), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1005), .ZN(new_n1304));
  OAI21_X1  g1104(.A(G390), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G396), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1305), .A2(new_n1290), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1307), .B1(new_n1305), .B2(new_n1290), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(G378), .B(new_n1257), .C1(new_n1262), .C2(new_n1265), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1231), .A2(new_n1264), .A3(new_n1268), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n828), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1232), .A2(new_n1256), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1294), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1298), .B1(new_n1311), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1267), .A2(KEYINPUT60), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1199), .A2(new_n1319), .A3(new_n1192), .A4(new_n1200), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1201), .A2(new_n1108), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1323), .A2(G384), .A3(new_n1285), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G384), .B1(new_n1323), .B2(new_n1285), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1317), .A2(KEYINPUT62), .A3(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1317), .B2(new_n1327), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1328), .A2(new_n1330), .A3(KEYINPUT126), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1317), .A2(new_n1327), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1329), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(KEYINPUT126), .A3(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1311), .A2(new_n1316), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1297), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1298), .A2(G2897), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1323), .A2(new_n1285), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n881), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1341), .A2(G2897), .A3(new_n1298), .A4(new_n1324), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1335), .B1(new_n1337), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1334), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1310), .B1(new_n1331), .B2(new_n1345), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1343), .A2(KEYINPUT123), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT123), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1339), .B2(new_n1342), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1317), .A2(KEYINPUT122), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1317), .A2(KEYINPUT122), .ZN(new_n1351));
  OAI22_X1  g1151(.A1(new_n1347), .A2(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(KEYINPUT63), .B1(new_n1317), .B2(new_n1327), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1353), .A2(new_n1310), .A3(KEYINPUT61), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1317), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1352), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1346), .A2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(G375), .A2(new_n1294), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1311), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT127), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1327), .A2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(KEYINPUT127), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1359), .A2(new_n1361), .A3(new_n1362), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1358), .A2(new_n1327), .A3(new_n1360), .A4(new_n1311), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  XOR2_X1   g1165(.A(new_n1365), .B(new_n1310), .Z(G402));
endmodule


