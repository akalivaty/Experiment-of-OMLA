//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215,
    new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(new_n440));
  INV_X1    g015(.A(new_n440), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n440), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n467), .A2(new_n474), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n467), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n474), .B2(G112), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT70), .Z(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n467), .A2(new_n488), .B1(new_n489), .B2(new_n463), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n463), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n490), .A2(G2105), .B1(G102), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n474), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n498), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G88), .ZN(new_n504));
  OAI21_X1  g079(.A(G543), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n510), .B(new_n511), .C1(new_n504), .C2(new_n503), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n498), .A2(new_n500), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT72), .A3(G62), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n505), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n530), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI211_X1 g108(.A(KEYINPUT73), .B(new_n532), .C1(new_n503), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n519), .A2(new_n509), .A3(G89), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT73), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n525), .B(new_n527), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n539));
  INV_X1    g114(.A(new_n527), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n532), .B1(new_n503), .B2(new_n533), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n540), .B1(new_n543), .B2(new_n534), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(new_n545), .A3(new_n525), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n539), .A2(new_n546), .ZN(G168));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  INV_X1    g123(.A(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n503), .A2(new_n548), .B1(new_n505), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n553), .B2(G651), .ZN(G171));
  NAND3_X1  g129(.A1(new_n519), .A2(new_n509), .A3(G81), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT76), .B(G43), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n505), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n519), .A2(G56), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT77), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n560), .B1(new_n515), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n505), .A2(new_n556), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n555), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT78), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G188));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n509), .A2(new_n579), .A3(G53), .A4(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n498), .A2(new_n500), .A3(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n578), .A2(new_n580), .B1(new_n583), .B2(G651), .ZN(new_n584));
  INV_X1    g159(.A(new_n503), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G91), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  NOR2_X1   g163(.A1(new_n538), .A2(KEYINPUT74), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n545), .B1(new_n544), .B2(new_n525), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(G286));
  NAND2_X1  g166(.A1(new_n585), .A2(G87), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n526), .A2(G49), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  AOI22_X1  g170(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT79), .B1(new_n596), .B2(new_n558), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n498), .A2(new_n500), .A3(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n600), .A2(new_n601), .A3(G651), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n597), .A2(new_n602), .B1(G86), .B2(new_n585), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n526), .A2(G48), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT80), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n585), .A2(G86), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n601), .B1(new_n600), .B2(G651), .ZN(new_n607));
  AOI211_X1 g182(.A(KEYINPUT79), .B(new_n558), .C1(new_n598), .C2(new_n599), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n604), .B(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n605), .A2(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT81), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  INV_X1    g190(.A(G85), .ZN(new_n616));
  INV_X1    g191(.A(G47), .ZN(new_n617));
  OAI22_X1  g192(.A1(new_n503), .A2(new_n616), .B1(new_n505), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(G290));
  AND3_X1   g195(.A1(new_n498), .A2(new_n500), .A3(G66), .ZN(new_n621));
  INV_X1    g196(.A(G79), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT83), .B1(new_n622), .B2(new_n497), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n624), .A2(G79), .A3(G543), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(G651), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G92), .ZN(new_n628));
  NOR2_X1   g203(.A1(KEYINPUT82), .A2(KEYINPUT10), .ZN(new_n629));
  AND2_X1   g204(.A1(KEYINPUT82), .A2(KEYINPUT10), .ZN(new_n630));
  OAI22_X1  g205(.A1(new_n503), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n526), .A2(G54), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n630), .A2(new_n629), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n519), .A2(new_n633), .A3(new_n509), .A4(G92), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n627), .A2(new_n631), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G171), .B2(new_n636), .ZN(G284));
  OAI21_X1  g213(.A(new_n637), .B1(G171), .B2(new_n636), .ZN(G321));
  NAND2_X1  g214(.A1(G299), .A2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G297));
  XNOR2_X1  g216(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g217(.A(new_n635), .ZN(new_n643));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(G860), .ZN(G148));
  INV_X1    g220(.A(new_n569), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(new_n636), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n635), .A2(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n636), .B2(new_n648), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g225(.A1(new_n464), .A2(new_n466), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n491), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT12), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n479), .A2(G123), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  OAI21_X1  g232(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n661), .C1(G111), .C2(new_n474), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n481), .A2(G135), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(G2096), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n655), .A2(new_n665), .ZN(G156));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2427), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2430), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT15), .B(G2435), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT14), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2451), .B(G2454), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2443), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2446), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n668), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n675), .A2(new_n678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n667), .A3(new_n679), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n682), .A2(G14), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n682), .A2(new_n684), .A3(KEYINPUT88), .A4(G14), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(G401));
  XOR2_X1   g264(.A(G2072), .B(G2078), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XNOR2_X1  g266(.A(G2084), .B(G2090), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2067), .B(G2678), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n697), .A2(KEYINPUT18), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(KEYINPUT18), .ZN(new_n699));
  OAI21_X1  g274(.A(KEYINPUT17), .B1(new_n693), .B2(new_n694), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n691), .B(new_n700), .Z(new_n701));
  OAI22_X1  g276(.A1(new_n698), .A2(new_n699), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G2100), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT91), .B(G2096), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(G2100), .ZN(new_n706));
  INV_X1    g281(.A(new_n704), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(G227));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1961), .B(G1966), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  XOR2_X1   g287(.A(G1956), .B(G2474), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1971), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT19), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n712), .A2(new_n713), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n719), .A2(new_n716), .A3(new_n714), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n714), .A2(new_n710), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(new_n718), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n717), .B(new_n720), .C1(new_n722), .C2(new_n716), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1991), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1981), .ZN(new_n726));
  XNOR2_X1  g301(.A(G1986), .B(G1996), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n724), .B(new_n728), .ZN(G229));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n643), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G4), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1348), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G35), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G162), .B2(new_n735), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2090), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n569), .A2(new_n730), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n730), .B2(G19), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT97), .B(G1341), .ZN(new_n742));
  AOI22_X1  g317(.A1(G1348), .A2(new_n733), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n739), .B(new_n743), .C1(new_n742), .C2(new_n741), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n745));
  INV_X1    g320(.A(G26), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G29), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n479), .A2(G128), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT98), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n481), .A2(G140), .ZN(new_n751));
  NOR2_X1   g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n745), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2067), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(G2067), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n578), .A2(new_n580), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n583), .A2(G651), .ZN(new_n760));
  AND3_X1   g335(.A1(new_n759), .A2(new_n586), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT23), .B1(new_n761), .B2(new_n730), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n730), .A2(G20), .ZN(new_n763));
  MUX2_X1   g338(.A(KEYINPUT23), .B(new_n762), .S(new_n763), .Z(new_n764));
  INV_X1    g339(.A(G1956), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n757), .A2(new_n758), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n738), .A2(G2090), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n744), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(G29), .A2(G32), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n479), .A2(G129), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT100), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n491), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n735), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n491), .A2(G103), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n481), .A2(G139), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n651), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n781), .B(new_n782), .C1(new_n474), .C2(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G33), .B(new_n784), .S(G29), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n777), .A2(new_n779), .B1(new_n785), .B2(G2072), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n735), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n735), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G2078), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n789), .C1(new_n777), .C2(new_n779), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT24), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n735), .B1(new_n791), .B2(G34), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n791), .A2(G34), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n477), .B2(new_n735), .ZN(new_n798));
  INV_X1    g373(.A(G2084), .ZN(new_n799));
  NOR2_X1   g374(.A1(G5), .A2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G171), .B2(G16), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n798), .A2(new_n799), .B1(G1961), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n799), .B2(new_n798), .ZN(new_n803));
  INV_X1    g378(.A(G28), .ZN(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n804), .B2(KEYINPUT30), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT30), .B2(new_n804), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n664), .B2(new_n735), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G2078), .B2(new_n788), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G1961), .B2(new_n801), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n785), .A2(G2072), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n790), .A2(new_n803), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G286), .A2(new_n730), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G1966), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT31), .B(G11), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n811), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n811), .A2(new_n818), .A3(new_n822), .A4(new_n819), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n769), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n603), .A2(KEYINPUT80), .A3(new_n604), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n609), .A2(new_n610), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n730), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(G6), .A2(G16), .ZN(new_n828));
  OR3_X1    g403(.A1(new_n827), .A2(KEYINPUT32), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT32), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G1981), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n730), .A2(G23), .ZN(new_n834));
  INV_X1    g409(.A(G288), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n730), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT33), .B(G1976), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n829), .A2(G1981), .A3(new_n830), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n730), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n730), .ZN(new_n842));
  INV_X1    g417(.A(G1971), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n833), .A2(new_n839), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT34), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(G119), .A2(new_n479), .B1(new_n481), .B2(G131), .ZN(new_n848));
  OR2_X1    g423(.A1(G95), .A2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n463), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .C1(G107), .C2(new_n474), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  MUX2_X1   g428(.A(G25), .B(new_n853), .S(G29), .Z(new_n854));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G1991), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT94), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n854), .B(new_n856), .Z(new_n857));
  NOR2_X1   g432(.A1(G16), .A2(G24), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT95), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(G16), .ZN(new_n860));
  INV_X1    g435(.A(G1986), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n847), .A2(new_n857), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT36), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n847), .A2(new_n865), .A3(new_n857), .A4(new_n862), .ZN(new_n866));
  AOI211_X1 g441(.A(new_n734), .B(new_n824), .C1(new_n864), .C2(new_n866), .ZN(G311));
  AOI21_X1  g442(.A(new_n824), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(G1348), .B2(new_n733), .ZN(G150));
  NAND3_X1  g444(.A1(new_n519), .A2(new_n509), .A3(G93), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n509), .A2(G55), .A3(G543), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT104), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT104), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(new_n558), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G860), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(KEYINPUT37), .Z(new_n880));
  AOI22_X1  g455(.A1(new_n875), .A2(new_n877), .B1(new_n562), .B2(new_n568), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n565), .A2(new_n555), .A3(new_n567), .ZN(new_n882));
  INV_X1    g457(.A(new_n874), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n882), .B(new_n877), .C1(new_n883), .C2(new_n872), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n635), .A2(new_n644), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT39), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n888), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n880), .B1(new_n891), .B2(G860), .ZN(G145));
  NAND2_X1  g467(.A1(new_n479), .A2(G130), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n481), .A2(G142), .ZN(new_n894));
  NOR2_X1   g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n664), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n486), .B(G160), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n776), .B(new_n853), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n486), .B(new_n477), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n898), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n754), .B(G164), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n784), .B(new_n653), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n904), .A3(new_n898), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n913), .B2(new_n905), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g492(.A1(new_n513), .A2(new_n522), .A3(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(G303), .A2(new_n835), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n919), .C1(new_n605), .C2(new_n611), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n513), .A2(new_n522), .A3(G288), .ZN(new_n921));
  AOI21_X1  g496(.A(G288), .B1(new_n513), .B2(new_n522), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n826), .B(new_n825), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n920), .A2(new_n923), .A3(new_n619), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n619), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AND4_X1   g503(.A1(KEYINPUT105), .A2(new_n635), .A3(new_n586), .A4(new_n584), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT105), .B1(new_n761), .B2(new_n635), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n643), .A2(G299), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n929), .B2(new_n930), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n643), .B2(G299), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n761), .A2(KEYINPUT105), .A3(new_n635), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT106), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n932), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n886), .B(new_n648), .ZN(new_n945));
  MUX2_X1   g520(.A(new_n933), .B(new_n944), .S(new_n945), .Z(new_n946));
  AND2_X1   g521(.A1(new_n928), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n928), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n878), .A2(new_n636), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(G295));
  XOR2_X1   g526(.A(G295), .B(KEYINPUT107), .Z(G331));
  NAND3_X1  g527(.A1(new_n539), .A2(new_n546), .A3(G171), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G171), .B1(new_n539), .B2(new_n546), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n954), .A2(new_n955), .B1(new_n885), .B2(new_n881), .ZN(new_n956));
  OAI21_X1  g531(.A(G301), .B1(new_n589), .B2(new_n590), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n886), .A3(new_n953), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n944), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n957), .A2(new_n886), .A3(KEYINPUT108), .A4(new_n953), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n962), .A2(new_n933), .A3(new_n956), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n960), .A2(new_n926), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n915), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n956), .A3(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n940), .A2(KEYINPUT41), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n931), .A2(new_n941), .A3(new_n932), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n956), .A2(new_n933), .A3(new_n958), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n924), .B2(new_n925), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n920), .A2(new_n923), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G290), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n920), .A2(new_n923), .A3(new_n619), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n966), .A2(new_n981), .A3(KEYINPUT43), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n965), .A2(new_n915), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n979), .B1(new_n960), .B2(new_n964), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT44), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n960), .A2(new_n964), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n983), .B1(new_n966), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n979), .B1(new_n970), .B2(new_n971), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n984), .A2(new_n993), .A3(KEYINPUT43), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n989), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n988), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n989), .B1(new_n982), .B2(new_n986), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n966), .A2(new_n981), .A3(new_n983), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT43), .B1(new_n984), .B2(new_n985), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT44), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(G397));
  XNOR2_X1  g578(.A(KEYINPUT111), .B(G1384), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n492), .B2(new_n494), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT112), .B(G40), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n476), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT126), .ZN(new_n1014));
  XOR2_X1   g589(.A(new_n754), .B(G2067), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1016), .B2(new_n776), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT125), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  NAND3_X1  g596(.A1(new_n1009), .A2(new_n861), .A3(new_n619), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT48), .Z(new_n1023));
  XNOR2_X1  g598(.A(new_n776), .B(G1996), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n853), .A2(new_n856), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n853), .A2(new_n856), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1023), .B1(new_n1029), .B2(new_n1009), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1009), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n754), .A2(G2067), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1021), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n476), .A2(new_n1007), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n492), .B2(new_n494), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1976), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(G288), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n832), .B1(new_n603), .B2(new_n604), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n609), .A2(G1981), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  OR3_X1    g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(G288), .B2(new_n1042), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1041), .B(new_n1051), .C1(new_n1042), .C2(G288), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n491), .A2(G102), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n489), .A2(new_n463), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n651), .B2(G126), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1060), .B2(new_n474), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT4), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n493), .B(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1055), .B(new_n1057), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1037), .A2(KEYINPUT115), .A3(new_n1057), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT116), .B(G2090), .Z(new_n1069));
  INV_X1    g644(.A(new_n1037), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT50), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1068), .A2(new_n1036), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1008), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1004), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT45), .B(new_n1077), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1005), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1036), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n843), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1073), .A2(new_n1076), .A3(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1087), .A2(G8), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G303), .A2(G8), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1089), .B(KEYINPUT55), .Z(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT118), .B(new_n1054), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1068), .A2(new_n799), .A3(new_n1036), .A4(new_n1071), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1037), .A2(KEYINPUT45), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n817), .B1(new_n1094), .B2(new_n1083), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(G8), .A3(G168), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1090), .B1(new_n1087), .B2(G8), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1053), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT63), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1054), .A2(KEYINPUT63), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1050), .A2(new_n1042), .A3(new_n835), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(G1981), .B2(new_n609), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1104), .A2(new_n1105), .B1(new_n1041), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n761), .B(KEYINPUT57), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT119), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1036), .B1(new_n1070), .B2(KEYINPUT50), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n765), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1082), .A2(new_n1084), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1110), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n635), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1038), .A2(G2067), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1068), .A2(new_n1036), .A3(new_n1071), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(G1348), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT60), .B(new_n1122), .C1(new_n1123), .C2(G1348), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n635), .A2(KEYINPUT122), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1068), .A2(new_n1036), .A3(new_n1071), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1121), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n635), .A2(KEYINPUT122), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n1133), .A4(new_n1127), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1082), .A2(new_n1084), .A3(new_n1010), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1038), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n569), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1144), .A3(new_n569), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(KEYINPUT59), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1118), .A2(KEYINPUT121), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1114), .A2(new_n1116), .A3(new_n1148), .A4(new_n1110), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1137), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1144), .B1(new_n1141), .B2(new_n569), .ZN(new_n1152));
  AOI211_X1 g727(.A(KEYINPUT120), .B(new_n646), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1110), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1119), .A2(new_n1155), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1154), .A2(KEYINPUT59), .B1(new_n1156), .B2(KEYINPUT61), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1125), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1159));
  INV_X1    g734(.A(G2078), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1082), .A2(new_n1084), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(G1961), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1130), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  INV_X1    g741(.A(new_n476), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1006), .A2(new_n1166), .A3(G40), .A4(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(G40), .B(new_n1167), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT124), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1162), .A2(G2078), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1168), .A2(new_n1170), .A3(new_n1082), .A4(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1163), .A2(new_n1165), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(G171), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1162), .A2(new_n1161), .B1(new_n1130), .B2(new_n1164), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1084), .A2(new_n1093), .A3(new_n1171), .ZN(new_n1176));
  AOI21_X1  g751(.A(G301), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1159), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1173), .A2(G171), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(G301), .A3(new_n1176), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(KEYINPUT54), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1092), .A2(G168), .A3(new_n1095), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(G8), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT51), .ZN(new_n1184));
  AOI21_X1  g759(.A(G168), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT51), .ZN(new_n1186));
  OAI211_X1 g761(.A(G8), .B(new_n1182), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1178), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1158), .A2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1097), .A2(KEYINPUT63), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1184), .A2(new_n1187), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1191), .B1(new_n1195), .B2(new_n1177), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1190), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1069), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1040), .B1(new_n1086), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1054), .B1(new_n1090), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1104), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1109), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1029), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n619), .B(G1986), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1031), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1035), .B1(new_n1203), .B2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  AOI22_X1  g782(.A1(new_n687), .A2(new_n688), .B1(new_n705), .B2(new_n708), .ZN(new_n1209));
  AND2_X1   g783(.A1(new_n1209), .A2(new_n916), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n999), .A2(new_n1000), .ZN(new_n1211));
  NOR2_X1   g785(.A1(G229), .A2(new_n460), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(G225));
  NAND2_X1  g787(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1214));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n1210), .A2(new_n1211), .A3(new_n1215), .A4(new_n1212), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1214), .A2(new_n1216), .ZN(G308));
endmodule


