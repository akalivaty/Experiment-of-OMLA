//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G97), .A2(G257), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G87), .A2(G250), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT69), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n212), .A2(new_n213), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n214), .B(new_n215), .C1(G77), .C2(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT70), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT71), .Z(new_n226));
  OR2_X1    g0026(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n227), .A2(G50), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT67), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT68), .Z(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n208), .A2(G13), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT0), .Z(new_n237));
  AND2_X1   g0037(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n238));
  NOR4_X1   g0038(.A1(new_n226), .A2(new_n234), .A3(new_n237), .A4(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT72), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT73), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT73), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G97), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n233), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(G33), .ZN(new_n266));
  AND4_X1   g0066(.A1(G97), .A2(new_n261), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT7), .B1(new_n270), .B2(new_n232), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT7), .ZN(new_n272));
  NOR4_X1   g0072(.A1(new_n268), .A2(new_n269), .A3(new_n272), .A4(G20), .ZN(new_n273));
  OAI21_X1  g0073(.A(G107), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT6), .ZN(new_n275));
  INV_X1    g0075(.A(G97), .ZN(new_n276));
  INV_X1    g0076(.A(G107), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G97), .A2(G107), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(KEYINPUT6), .A3(G97), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G20), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G77), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n274), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI211_X1 g0086(.A(new_n262), .B(new_n267), .C1(new_n286), .C2(new_n264), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  OAI211_X1 g0089(.A(G1), .B(G13), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n260), .A2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT84), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(new_n289), .A3(KEYINPUT5), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT5), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(KEYINPUT84), .B2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(G257), .B(new_n290), .C1(new_n291), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  INV_X1    g0098(.A(G45), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n257), .B2(new_n259), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n298), .A2(G274), .A3(new_n290), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  OAI211_X1 g0104(.A(G244), .B(new_n304), .C1(new_n268), .C2(new_n269), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT4), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT3), .B(G33), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(KEYINPUT4), .A3(G244), .A4(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G283), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(G250), .A3(G1698), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n302), .B1(new_n303), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G190), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n303), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT83), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT83), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n317), .A3(new_n303), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n302), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n287), .B(new_n314), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  OAI211_X1 g0121(.A(G257), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n322));
  OAI211_X1 g0122(.A(G250), .B(new_n304), .C1(new_n268), .C2(new_n269), .ZN(new_n323));
  INV_X1    g0123(.A(G294), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n322), .B(new_n323), .C1(new_n288), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n303), .ZN(new_n326));
  OAI211_X1 g0126(.A(G264), .B(new_n290), .C1(new_n291), .C2(new_n296), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n301), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n320), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n326), .A2(new_n330), .A3(new_n301), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n261), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT25), .A3(new_n277), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT25), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n261), .B2(G107), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(new_n336), .B1(new_n337), .B2(G107), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n232), .B(G87), .C1(new_n268), .C2(new_n269), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT87), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT22), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n308), .A2(new_n232), .A3(G87), .A4(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n232), .A2(G33), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G116), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n232), .A2(G107), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT23), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n343), .A2(new_n344), .B1(G116), .B2(new_n347), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(new_n350), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n353), .A2(new_n356), .B1(KEYINPUT88), .B2(KEYINPUT24), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n332), .B(new_n338), .C1(new_n357), .C2(new_n265), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n297), .A2(new_n301), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n312), .A2(new_n317), .A3(new_n303), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n317), .B1(new_n312), .B2(new_n303), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n315), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n267), .ZN(new_n367));
  INV_X1    g0167(.A(new_n262), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n272), .B1(new_n308), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n277), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n285), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n232), .B1(new_n280), .B2(new_n281), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n367), .B(new_n368), .C1(new_n374), .C2(new_n265), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n363), .A2(new_n366), .A3(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n321), .A2(new_n358), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G41), .A2(G45), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n256), .A3(G274), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT73), .B(G1), .ZN(new_n381));
  OAI211_X1 g0181(.A(G238), .B(new_n290), .C1(new_n381), .C2(new_n378), .ZN(new_n382));
  OR2_X1    g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  INV_X1    g0184(.A(G232), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n217), .A2(new_n304), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(new_n387), .B1(G33), .B2(G97), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n380), .B(new_n382), .C1(new_n388), .C2(new_n290), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT13), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n387), .B1(G232), .B2(new_n304), .C1(new_n268), .C2(new_n269), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n303), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n380), .A4(new_n382), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n389), .A2(new_n398), .A3(KEYINPUT13), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G179), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n396), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G169), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT14), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n365), .B1(new_n390), .B2(new_n396), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n333), .A2(new_n218), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT12), .ZN(new_n410));
  OR3_X1    g0210(.A1(new_n381), .A2(KEYINPUT76), .A3(new_n232), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT76), .B1(new_n381), .B2(new_n232), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n265), .A4(new_n261), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G68), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n284), .A2(G50), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(new_n232), .B2(G68), .C1(new_n203), .C2(new_n346), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n264), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT11), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n410), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n408), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n400), .A2(G190), .ZN(new_n422));
  INV_X1    g0222(.A(new_n420), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n402), .A2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(KEYINPUT80), .A3(new_n425), .ZN(new_n429));
  INV_X1    g0229(.A(new_n380), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n308), .A2(G238), .A3(G1698), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n308), .A2(G232), .A3(new_n304), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n277), .C2(new_n308), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(new_n303), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT77), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n303), .B1(new_n260), .B2(new_n379), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G244), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n435), .B1(new_n434), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n359), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n440), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(new_n365), .A3(new_n438), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n414), .A2(G77), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n333), .A2(new_n203), .ZN(new_n445));
  XOR2_X1   g0245(.A(KEYINPUT8), .B(G58), .Z(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT15), .B(G87), .Z(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n346), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n264), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n441), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n428), .A2(new_n429), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n333), .A2(new_n202), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n232), .B1(new_n201), .B2(new_n202), .ZN(new_n456));
  INV_X1    g0256(.A(G150), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n457), .A2(G20), .A3(G33), .ZN(new_n458));
  INV_X1    g0258(.A(G58), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT74), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT75), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G58), .ZN(new_n462));
  OAI211_X1 g0262(.A(KEYINPUT8), .B(new_n460), .C1(new_n462), .C2(KEYINPUT74), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n462), .A2(KEYINPUT8), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI211_X1 g0265(.A(new_n456), .B(new_n458), .C1(new_n465), .C2(new_n347), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n455), .B1(new_n413), .B2(new_n202), .C1(new_n466), .C2(new_n265), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT9), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G222), .A2(G1698), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n304), .A2(G223), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n308), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n473), .B(new_n303), .C1(G77), .C2(new_n308), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n290), .B1(new_n381), .B2(new_n378), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(new_n380), .C1(new_n217), .C2(new_n475), .ZN(new_n476));
  XOR2_X1   g0276(.A(KEYINPUT78), .B(G200), .Z(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n476), .A2(new_n330), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n469), .A2(new_n470), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT10), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n476), .A2(G179), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n365), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n467), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n475), .A2(new_n385), .ZN(new_n486));
  OR2_X1    g0286(.A1(G223), .A2(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n217), .A2(G1698), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n268), .C2(new_n269), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G87), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n290), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR4_X1   g0291(.A1(new_n486), .A2(new_n491), .A3(G179), .A4(new_n430), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n490), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n430), .B1(new_n493), .B2(new_n303), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n436), .A2(G232), .ZN(new_n495));
  AOI21_X1  g0295(.A(G169), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT82), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n359), .A3(new_n495), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n486), .A2(new_n491), .A3(new_n430), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n498), .B(new_n499), .C1(new_n500), .C2(G169), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n284), .A2(G159), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT74), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G58), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n460), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n201), .B1(new_n506), .B2(G68), .ZN(new_n507));
  OAI211_X1 g0307(.A(KEYINPUT81), .B(new_n503), .C1(new_n507), .C2(new_n232), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT16), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n503), .B1(new_n507), .B2(new_n232), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n218), .B1(new_n369), .B2(new_n370), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n201), .ZN(new_n513));
  XNOR2_X1  g0313(.A(KEYINPUT74), .B(G58), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n218), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G20), .B1(G159), .B2(new_n284), .ZN(new_n516));
  OAI21_X1  g0316(.A(G68), .B1(new_n271), .B2(new_n273), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n516), .B(new_n517), .C1(KEYINPUT81), .C2(KEYINPUT16), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n512), .A2(new_n518), .A3(new_n264), .ZN(new_n519));
  INV_X1    g0319(.A(new_n465), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n261), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n414), .B2(new_n520), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT18), .B1(new_n502), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n502), .A2(KEYINPUT18), .A3(new_n523), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n494), .A2(new_n330), .A3(new_n495), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n500), .B2(G200), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n519), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT17), .ZN(new_n531));
  OAI21_X1  g0331(.A(G190), .B1(new_n439), .B2(new_n440), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n442), .A2(new_n477), .A3(new_n438), .ZN(new_n533));
  INV_X1    g0333(.A(new_n452), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n527), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n454), .A2(new_n485), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n261), .A2(new_n266), .A3(new_n265), .A4(G116), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n333), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(G20), .B1(G33), .B2(G283), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n288), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT86), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT86), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n263), .A2(new_n233), .B1(G20), .B2(new_n540), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT86), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT86), .B1(new_n542), .B2(new_n543), .ZN(new_n552));
  OAI211_X1 g0352(.A(KEYINPUT20), .B(new_n549), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n539), .B(new_n541), .C1(new_n550), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G264), .B(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(new_n304), .C1(new_n268), .C2(new_n269), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n383), .A2(G303), .A3(new_n384), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n303), .ZN(new_n561));
  OAI211_X1 g0361(.A(G270), .B(new_n290), .C1(new_n291), .C2(new_n296), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n301), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G169), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n538), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n563), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G190), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n555), .A2(G179), .A3(new_n566), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n563), .A2(G169), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(KEYINPUT21), .A3(new_n555), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n219), .A2(new_n304), .ZN(new_n574));
  INV_X1    g0374(.A(G244), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G1698), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n576), .C1(new_n268), .C2(new_n269), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n303), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n300), .A2(G274), .A3(new_n290), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n291), .A2(G250), .A3(new_n290), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n359), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n583), .B(KEYINPUT85), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n365), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n232), .B1(new_n392), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n279), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n232), .B(G68), .C1(new_n268), .C2(new_n269), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n346), .B2(new_n276), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n264), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n381), .A2(new_n232), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n449), .A2(new_n596), .A3(G13), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n261), .A2(new_n266), .A3(new_n265), .A4(new_n448), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n586), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n585), .A2(new_n330), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n261), .A2(new_n266), .A3(new_n265), .A4(G87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n585), .A2(new_n477), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n584), .A2(new_n600), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n573), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n338), .B1(new_n357), .B2(new_n265), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n328), .A2(new_n365), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n303), .B1(new_n298), .B2(new_n300), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(G264), .B1(new_n325), .B2(new_n303), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n359), .A3(new_n301), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n377), .A2(new_n537), .A3(new_n608), .A4(new_n614), .ZN(G372));
  AND3_X1   g0415(.A1(new_n586), .A2(new_n599), .A3(new_n583), .ZN(new_n616));
  INV_X1    g0416(.A(new_n477), .ZN(new_n617));
  INV_X1    g0417(.A(new_n581), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n290), .B1(new_n577), .B2(new_n578), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n582), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT89), .B1(new_n621), .B2(new_n603), .ZN(new_n622));
  INV_X1    g0422(.A(new_n601), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n604), .A2(new_n605), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n376), .A2(new_n321), .A3(new_n358), .A4(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n571), .A2(KEYINPUT21), .A3(new_n555), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT21), .B1(new_n571), .B2(new_n555), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n555), .A2(G179), .A3(new_n566), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n614), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n616), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT26), .B1(new_n607), .B2(new_n376), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n603), .B1(new_n585), .B2(new_n477), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n601), .B1(new_n635), .B2(new_n624), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n616), .B1(new_n636), .B2(new_n622), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n376), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n363), .A2(new_n375), .A3(new_n366), .A4(KEYINPUT90), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n633), .B(new_n634), .C1(KEYINPUT26), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n537), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n484), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n400), .A2(G179), .B1(new_n406), .B2(new_n405), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n423), .B1(new_n645), .B2(new_n404), .ZN(new_n646));
  INV_X1    g0446(.A(new_n453), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n425), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT17), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n530), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n527), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n644), .B1(new_n651), .B2(new_n481), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n643), .A2(new_n652), .ZN(G369));
  NAND2_X1  g0453(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n351), .A2(new_n352), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n355), .B1(new_n354), .B2(new_n350), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n264), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n658), .A2(new_n338), .B1(new_n365), .B2(new_n328), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n232), .A2(G13), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n381), .A2(KEYINPUT91), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  INV_X1    g0462(.A(new_n660), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n260), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n661), .A2(new_n664), .A3(KEYINPUT27), .ZN(new_n665));
  INV_X1    g0465(.A(G213), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT27), .B1(new_n661), .B2(new_n664), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT92), .B(KEYINPUT27), .C1(new_n661), .C2(new_n664), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n609), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n659), .A2(new_n613), .B1(new_n675), .B2(new_n358), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n614), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT94), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n614), .ZN(new_n679));
  INV_X1    g0479(.A(new_n674), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n358), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n614), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n631), .B(new_n569), .C1(new_n556), .C2(new_n680), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n565), .A2(new_n570), .A3(new_n572), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n555), .A3(new_n674), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT93), .B(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n631), .A2(new_n674), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n678), .A2(new_n685), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT95), .A3(new_n681), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT95), .B1(new_n698), .B2(new_n681), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n700), .B2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n235), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n590), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT96), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n230), .B2(new_n704), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(KEYINPUT96), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT98), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n607), .A2(new_n376), .A3(KEYINPUT26), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n633), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n716), .B2(new_n680), .ZN(new_n717));
  AOI211_X1 g0517(.A(KEYINPUT98), .B(new_n674), .C1(new_n633), .C2(new_n715), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT29), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n642), .A2(new_n680), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n608), .A2(new_n377), .A3(new_n614), .A4(new_n680), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT97), .B(KEYINPUT31), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n359), .A3(new_n328), .A4(new_n563), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n562), .A2(new_n301), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n612), .A3(G179), .A4(new_n561), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(new_n360), .A3(new_n315), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n561), .A2(new_n562), .A3(new_n301), .A4(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n326), .A2(new_n327), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n313), .A3(KEYINPUT30), .A4(new_n729), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n674), .B(new_n726), .C1(new_n730), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n319), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n328), .A3(new_n585), .A4(new_n563), .ZN(new_n743));
  INV_X1    g0543(.A(new_n740), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n680), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n741), .B1(new_n745), .B2(KEYINPUT31), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n693), .B1(new_n725), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n723), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n712), .B1(new_n749), .B2(G1), .ZN(G364));
  INV_X1    g0550(.A(new_n695), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n692), .A2(new_n694), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n256), .B1(new_n663), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n704), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n251), .A2(G45), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n703), .A2(new_n308), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(new_n231), .C2(G45), .ZN(new_n760));
  NAND3_X1  g0560(.A1(G355), .A2(new_n235), .A3(new_n308), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n761), .C1(G116), .C2(new_n235), .ZN(new_n762));
  INV_X1    g0562(.A(G13), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n288), .A3(KEYINPUT99), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT99), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G13), .B2(G33), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n233), .B1(G20), .B2(new_n365), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT100), .Z(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n232), .B1(new_n774), .B2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n276), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n232), .A2(new_n330), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n359), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n232), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n779), .A2(new_n514), .B1(new_n781), .B2(new_n203), .ZN(new_n782));
  NAND3_X1  g0582(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n776), .B(new_n782), .C1(G68), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n774), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n477), .A2(new_n359), .A3(new_n780), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(KEYINPUT32), .B1(new_n790), .B2(new_n277), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n477), .A2(new_n359), .A3(new_n777), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n589), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n783), .A2(new_n330), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G50), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n270), .B1(new_n789), .B2(KEYINPUT32), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n785), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n790), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n779), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n308), .B(new_n801), .C1(G322), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n786), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G329), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n781), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n784), .ZN(new_n808));
  INV_X1    g0608(.A(G317), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n809), .A2(KEYINPUT33), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(KEYINPUT33), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n807), .B(new_n812), .C1(G326), .C2(new_n795), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n803), .A2(new_n805), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n775), .A2(new_n324), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n798), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n762), .A2(new_n773), .B1(new_n770), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n769), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n691), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n757), .B1(new_n756), .B2(new_n819), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n453), .A2(new_n674), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n535), .B1(new_n534), .B2(new_n680), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n453), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n720), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n616), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n689), .B1(new_n659), .B2(new_n613), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n321), .A2(new_n358), .A3(new_n626), .A4(new_n376), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n634), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n823), .B(new_n680), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(new_n747), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n756), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n824), .A2(new_n767), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n790), .A2(new_n589), .B1(new_n806), .B2(new_n786), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT102), .Z(new_n837));
  INV_X1    g0637(.A(new_n781), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G294), .A2(new_n802), .B1(new_n838), .B2(G116), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n776), .B1(new_n784), .B2(G283), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n308), .B1(new_n795), .B2(G303), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n837), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n792), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(G107), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n790), .A2(new_n218), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n802), .A2(G143), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G137), .A2(new_n795), .B1(new_n784), .B2(G150), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(new_n787), .C2(new_n781), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n846), .B1(new_n202), .B2(new_n792), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n270), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n853), .B2(new_n786), .ZN(new_n854));
  INV_X1    g0654(.A(new_n775), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n851), .B(new_n854), .C1(new_n506), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n770), .B1(new_n844), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n767), .A2(new_n770), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n203), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n835), .A2(new_n755), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n834), .A2(new_n860), .ZN(G384));
  INV_X1    g0661(.A(new_n672), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT16), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n264), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n522), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n502), .A2(KEYINPUT18), .A3(new_n523), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n524), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n862), .B(new_n866), .C1(new_n868), .C2(new_n650), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n502), .A2(new_n523), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n519), .A2(new_n522), .A3(new_n529), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n672), .B1(new_n519), .B2(new_n522), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n502), .A2(new_n523), .A3(KEYINPUT104), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n872), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n502), .A2(new_n866), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n866), .A2(new_n862), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n530), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n523), .A2(new_n862), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n870), .A2(new_n885), .A3(new_n530), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n878), .A2(KEYINPUT105), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT105), .B1(new_n878), .B2(new_n887), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n885), .B1(new_n527), .B2(new_n531), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n884), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT103), .B1(new_n646), .B2(new_n674), .ZN(new_n893));
  AND4_X1   g0693(.A1(KEYINPUT103), .A2(new_n408), .A3(new_n420), .A4(new_n674), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n680), .A2(new_n423), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n893), .A2(new_n894), .B1(new_n426), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n726), .ZN(new_n897));
  INV_X1    g0697(.A(new_n728), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n740), .B1(new_n898), .B2(new_n585), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n899), .B2(new_n680), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT31), .B(new_n674), .C1(new_n730), .C2(new_n740), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n724), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n823), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n896), .A4(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n878), .A2(new_n882), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n880), .B1(new_n527), .B2(new_n531), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n884), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n896), .A3(new_n903), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n537), .A2(new_n902), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n913), .B(new_n914), .Z(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n693), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n719), .A2(new_n537), .A3(new_n722), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n652), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n421), .A2(new_n674), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n884), .C1(new_n891), .C2(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n821), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n831), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n909), .A2(new_n928), .A3(new_n896), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n527), .A2(new_n862), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n920), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n426), .ZN(new_n934));
  INV_X1    g0734(.A(new_n895), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT103), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n421), .B2(new_n680), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n646), .A2(KEYINPUT103), .A3(new_n674), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n934), .A2(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n831), .B2(new_n927), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n930), .B1(new_n940), .B2(new_n909), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n923), .B1(new_n908), .B2(new_n884), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n869), .A2(new_n883), .A3(KEYINPUT38), .ZN(new_n943));
  INV_X1    g0743(.A(new_n890), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n878), .A2(new_n887), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT105), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n878), .A2(KEYINPUT105), .A3(new_n887), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n949), .B2(new_n905), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n942), .B1(new_n950), .B2(new_n923), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n941), .B(KEYINPUT106), .C1(new_n951), .C2(new_n922), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n933), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n919), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n260), .B2(new_n663), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n540), .B1(new_n282), .B2(KEYINPUT35), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n233), .A2(new_n232), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(KEYINPUT35), .C2(new_n282), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT36), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n230), .B(G77), .C1(new_n218), .C2(new_n514), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(G50), .B2(new_n218), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n961), .A2(new_n763), .A3(new_n381), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n955), .A2(new_n959), .A3(new_n962), .ZN(G367));
  OAI211_X1 g0763(.A(new_n321), .B(new_n376), .C1(new_n680), .C2(new_n287), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n376), .B2(new_n680), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT109), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT42), .B1(new_n967), .B2(new_n698), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n679), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n376), .ZN(new_n970));
  OAI211_X1 g0770(.A(KEYINPUT110), .B(new_n968), .C1(new_n970), .C2(new_n674), .ZN(new_n971));
  INV_X1    g0771(.A(new_n698), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT42), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n966), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT110), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n674), .B1(new_n969), .B2(new_n376), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n973), .B1(new_n972), .B2(new_n966), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n637), .B1(new_n604), .B2(new_n680), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT107), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n680), .A2(new_n604), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n980), .A2(new_n981), .B1(new_n616), .B2(new_n982), .ZN(new_n983));
  NOR4_X1   g0783(.A1(new_n680), .A2(new_n826), .A3(KEYINPUT107), .A4(new_n604), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n979), .A2(new_n987), .A3(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n991), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n971), .A2(new_n978), .A3(new_n993), .A4(new_n974), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n696), .A2(new_n967), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n704), .B(KEYINPUT41), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n966), .B1(new_n700), .B2(new_n701), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(KEYINPUT45), .B(new_n966), .C1(new_n700), .C2(new_n701), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n701), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1005), .A2(new_n699), .A3(new_n967), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1005), .A2(KEYINPUT44), .A3(new_n699), .A4(new_n967), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n696), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n751), .A2(new_n686), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n696), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n697), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n748), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1004), .A2(new_n1010), .A3(new_n696), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1013), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1020), .B2(new_n749), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n997), .B1(new_n1021), .B2(new_n754), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n772), .B1(new_n247), .B2(new_n759), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n448), .A2(new_n703), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n756), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n838), .A2(G50), .B1(G159), .B2(new_n784), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n308), .C1(new_n457), .C2(new_n779), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n795), .A2(G143), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n218), .B2(new_n775), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n843), .B2(new_n506), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1031), .B1(new_n203), .B2(new_n790), .C1(new_n1032), .C2(new_n786), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n808), .A2(new_n324), .B1(new_n779), .B2(new_n800), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G317), .B2(new_n804), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n308), .B1(new_n838), .B2(G283), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n790), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(G97), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n855), .A2(G107), .B1(G311), .B2(new_n795), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n792), .A2(new_n540), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT46), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1028), .A2(new_n1033), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT47), .Z(new_n1044));
  INV_X1    g0844(.A(new_n770), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1025), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT112), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n986), .B2(new_n818), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1022), .A2(new_n1048), .ZN(G387));
  INV_X1    g0849(.A(new_n1018), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1017), .A2(new_n748), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n704), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n756), .B1(new_n686), .B2(new_n769), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n446), .A2(new_n202), .ZN(new_n1054));
  XOR2_X1   g0854(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n706), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n759), .C1(new_n243), .C2(new_n299), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n308), .A2(new_n235), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(G107), .B2(new_n235), .C1(new_n706), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n773), .A2(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n779), .A2(new_n202), .B1(new_n781), .B2(new_n218), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n795), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1038), .B1(new_n787), .B2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n792), .A2(new_n203), .B1(new_n457), .B2(new_n786), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1063), .B(new_n1065), .C1(KEYINPUT114), .C2(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(KEYINPUT114), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n465), .A2(new_n784), .B1(new_n448), .B2(new_n855), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1067), .A2(new_n308), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G311), .A2(new_n784), .B1(new_n795), .B2(G322), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n800), .B2(new_n781), .C1(new_n809), .C2(new_n779), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT48), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n799), .B2(new_n775), .C1(new_n324), .C2(new_n792), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT49), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n804), .A2(G326), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1076), .B(new_n270), .C1(new_n790), .C2(new_n540), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n770), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1053), .A2(new_n1062), .A3(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1052), .B(new_n1080), .C1(new_n753), .C2(new_n1017), .ZN(G393));
  NAND3_X1  g0881(.A1(new_n1013), .A2(new_n754), .A3(new_n1019), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n756), .B1(new_n967), .B2(new_n769), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n772), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n759), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1084), .B1(new_n276), .B2(new_n235), .C1(new_n254), .C2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n802), .A2(G159), .B1(G150), .B2(new_n795), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT51), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n446), .B2(new_n838), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n218), .A2(new_n792), .B1(new_n790), .B2(new_n589), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n270), .B(new_n1090), .C1(G50), .C2(new_n784), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n855), .A2(G77), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n804), .A2(G143), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n802), .A2(G311), .B1(G317), .B2(new_n795), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT52), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n308), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n781), .A2(new_n324), .B1(new_n775), .B2(new_n540), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G303), .B2(new_n784), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT115), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n804), .A2(G322), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G107), .A2(new_n1037), .B1(new_n843), .B2(G283), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1094), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1083), .B(new_n1086), .C1(new_n1045), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1082), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n705), .B1(new_n1107), .B2(new_n1050), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n1108), .B2(new_n1020), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(G390));
  NAND3_X1  g0910(.A1(new_n537), .A2(G330), .A3(new_n902), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n917), .A2(new_n652), .A3(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n693), .B(new_n823), .C1(new_n725), .C2(new_n746), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n939), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT116), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n903), .A2(new_n1116), .A3(G330), .A4(new_n896), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n896), .A2(G330), .A3(new_n823), .A4(new_n902), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1113), .A2(new_n939), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n928), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1113), .A2(new_n939), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n641), .A2(KEYINPUT26), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n714), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n680), .B1(new_n1127), .B2(new_n829), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT98), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n716), .A2(new_n713), .A3(new_n680), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(new_n927), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n822), .A2(new_n453), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n903), .A2(G330), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n939), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1112), .B1(new_n1123), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n1132), .A3(new_n896), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n950), .A2(new_n921), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n924), .B(new_n925), .C1(new_n940), .C2(new_n921), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1124), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n704), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n1137), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT118), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n1149), .A3(new_n704), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n754), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n951), .A2(new_n767), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n756), .B1(new_n520), .B2(new_n858), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n843), .A2(G150), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT53), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT54), .B(G143), .Z(new_n1157));
  AOI22_X1  g0957(.A1(new_n838), .A2(new_n1157), .B1(G137), .B2(new_n784), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT119), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n795), .A2(G128), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n787), .C2(new_n775), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G50), .B2(new_n1037), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n804), .A2(G125), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n308), .A3(new_n1163), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1156), .B(new_n1164), .C1(G132), .C2(new_n802), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n793), .B1(G116), .B2(new_n802), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n799), .B2(new_n1064), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G294), .B2(new_n804), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n270), .B1(new_n808), .B2(new_n277), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G97), .B2(new_n838), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n846), .A3(new_n1092), .A4(new_n1170), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  OAI21_X1  g0972(.A(new_n770), .B1(new_n1165), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1153), .A2(new_n1154), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1152), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1152), .A2(KEYINPUT121), .A3(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1151), .A2(new_n1179), .ZN(G378));
  INV_X1    g0980(.A(new_n1112), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1145), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n904), .A2(new_n912), .A3(G330), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n953), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n862), .A2(new_n467), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n485), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT124), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n933), .A2(new_n952), .A3(new_n1183), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1190), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n933), .A2(new_n952), .A3(new_n1183), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1183), .B1(new_n933), .B2(new_n952), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1182), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1182), .A2(new_n1196), .A3(new_n1192), .A4(KEYINPUT57), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n704), .A3(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1192), .A3(new_n754), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n808), .A2(new_n276), .B1(new_n775), .B2(new_n218), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1037), .A2(new_n506), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n270), .C1(new_n799), .C2(new_n786), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G41), .B(new_n1205), .C1(G77), .C2(new_n843), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT123), .Z(new_n1207));
  AOI211_X1 g1007(.A(new_n1203), .B(new_n1207), .C1(new_n448), .C2(new_n838), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n277), .B2(new_n779), .C1(new_n540), .C2(new_n1064), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT58), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n843), .A2(new_n1157), .B1(G128), .B2(new_n802), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n795), .A2(G125), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n855), .A2(G150), .B1(G132), .B2(new_n784), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G137), .B2(new_n838), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n804), .C2(G124), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(new_n787), .C2(new_n790), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G50), .B1(new_n384), .B2(new_n289), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1210), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n770), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n858), .A2(new_n202), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1189), .A2(new_n768), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n755), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1202), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1201), .A2(new_n1226), .ZN(G375));
  INV_X1    g1027(.A(new_n1137), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1123), .A2(new_n1112), .A3(new_n1136), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n998), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n753), .B1(new_n1123), .B2(new_n1136), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n939), .A2(new_n767), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1157), .A2(new_n784), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1233), .B(new_n308), .C1(new_n202), .C2(new_n775), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G150), .A2(new_n838), .B1(new_n804), .B2(G128), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1204), .A2(new_n1235), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1032), .B2(new_n779), .C1(new_n787), .C2(new_n792), .ZN(new_n1237));
  AOI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(G132), .C2(new_n795), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n308), .B1(new_n784), .B2(G116), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n324), .B2(new_n1064), .C1(new_n449), .C2(new_n775), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G283), .A2(new_n802), .B1(new_n838), .B2(G107), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n203), .B2(new_n790), .C1(new_n800), .C2(new_n786), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1240), .B(new_n1242), .C1(G97), .C2(new_n843), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n770), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n858), .A2(new_n218), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1232), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1231), .B1(new_n755), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1230), .A2(new_n1247), .ZN(G381));
  XOR2_X1   g1048(.A(G375), .B(KEYINPUT125), .Z(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G378), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1022), .A2(new_n1048), .A3(new_n1109), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1251), .A2(G396), .A3(G393), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G381), .A2(G384), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(G407));
  AOI21_X1  g1054(.A(new_n666), .B1(new_n1250), .B2(new_n673), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(G407), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n1201), .A2(G378), .A3(new_n1226), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1202), .B(new_n1225), .C1(new_n1197), .C2(new_n999), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(new_n1179), .A3(new_n1151), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n666), .A2(G343), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1229), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1229), .A2(new_n1263), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n704), .A3(new_n1228), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1266), .B2(new_n1247), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(G384), .A3(new_n1247), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1260), .A2(new_n1262), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1269), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G2897), .B(new_n1261), .C1(new_n1275), .C2(new_n1267), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1261), .A2(G2897), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1268), .A2(new_n1269), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1274), .A2(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1260), .A2(new_n1283), .A3(new_n1262), .A4(new_n1271), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1273), .A2(new_n1281), .A3(new_n1282), .A4(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(G396), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1251), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1109), .B1(new_n1022), .B2(new_n1048), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(G390), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1251), .A3(new_n1286), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1285), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1279), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1261), .B(new_n1270), .C1(new_n1257), .C2(new_n1259), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT63), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1290), .A2(new_n1292), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT126), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1272), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1290), .A2(new_n1292), .A3(new_n1303), .A4(new_n1298), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1297), .A2(new_n1300), .A3(new_n1302), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1294), .A2(new_n1305), .ZN(G405));
  INV_X1    g1106(.A(new_n1257), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G378), .B1(new_n1201), .B2(new_n1226), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1293), .A2(new_n1309), .ZN(new_n1310));
  OAI211_X1 g1110(.A(new_n1290), .B(new_n1292), .C1(new_n1308), .C2(new_n1307), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1270), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1271), .A3(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G402));
endmodule


