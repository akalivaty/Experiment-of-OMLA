//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n192), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT11), .B1(new_n201), .B2(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G134), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(new_n201), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(G137), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT11), .A2(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n216), .B2(G137), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n201), .A3(G134), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT64), .A2(G137), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT64), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n210), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n200), .B1(new_n215), .B2(new_n225), .ZN(new_n226));
  AOI211_X1 g040(.A(KEYINPUT67), .B(new_n224), .C1(new_n212), .C2(new_n214), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n199), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n204), .A2(new_n209), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n212), .A2(new_n214), .B1(G131), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n190), .A2(new_n192), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n190), .A2(new_n192), .A3(new_n232), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n243), .A2(new_n247), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n215), .A2(new_n225), .A3(new_n199), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n233), .B2(new_n234), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n190), .A2(new_n192), .A3(new_n232), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n231), .A2(new_n232), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n190), .A2(new_n192), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT69), .B(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n251), .B(new_n252), .C1(new_n230), .C2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n238), .A2(new_n250), .B1(KEYINPUT72), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n262), .B(new_n252), .C1(new_n228), .C2(new_n237), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n188), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G101), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT30), .B1(new_n228), .B2(new_n237), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n229), .A2(G131), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n215), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n254), .A2(new_n258), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n251), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n277), .A2(new_n252), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n260), .A2(new_n274), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n276), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n224), .B1(new_n212), .B2(new_n214), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(new_n200), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n236), .B1(new_n292), .B2(new_n199), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n250), .B(new_n290), .C1(new_n293), .C2(KEYINPUT30), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n274), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT70), .B1(new_n260), .B2(new_n274), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n269), .A2(new_n275), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n187), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n283), .A2(new_n288), .A3(new_n276), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT31), .B1(new_n294), .B2(new_n297), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n274), .B1(new_n264), .B2(new_n268), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT74), .B(new_n300), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n302), .A2(new_n308), .A3(new_n311), .A4(new_n303), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n299), .A2(new_n301), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT32), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n260), .A2(KEYINPUT76), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n279), .A2(new_n280), .B1(new_n291), .B2(new_n199), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n252), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n260), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n268), .B1(new_n265), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n269), .A2(new_n321), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n275), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n294), .A2(new_n260), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n274), .ZN(new_n326));
  AOI21_X1  g140(.A(G902), .B1(new_n326), .B2(new_n321), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G472), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n310), .A2(new_n312), .A3(new_n314), .A4(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G122), .ZN(new_n333));
  INV_X1    g147(.A(G104), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n334), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G104), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(G107), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G101), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n335), .A2(new_n338), .A3(new_n342), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n345), .A3(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n250), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n250), .A2(KEYINPUT84), .A3(new_n344), .A4(new_n346), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n334), .A2(G107), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n337), .A2(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(G101), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n245), .B2(new_n246), .ZN(new_n357));
  OAI21_X1  g171(.A(G113), .B1(new_n240), .B2(KEYINPUT5), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(new_n249), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n350), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT85), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n349), .A2(new_n362), .A3(new_n350), .A4(new_n359), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n333), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT6), .ZN(new_n365));
  INV_X1    g179(.A(new_n333), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT6), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n198), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n371), .B(KEYINPUT88), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n235), .A2(G125), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n235), .A2(KEYINPUT86), .A3(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT87), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n372), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n372), .A2(new_n379), .A3(KEYINPUT89), .A4(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G224), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n369), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(KEYINPUT7), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n371), .B(KEYINPUT88), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n377), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n333), .B(KEYINPUT8), .Z(new_n396));
  NOR2_X1   g210(.A1(new_n243), .A2(new_n356), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n249), .B1(new_n397), .B2(new_n358), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n398), .B2(new_n355), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n249), .B1(new_n357), .B2(new_n358), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(new_n355), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n387), .B(KEYINPUT90), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n404));
  OAI221_X1 g218(.A(new_n402), .B1(new_n381), .B2(new_n404), .C1(new_n360), .C2(new_n366), .ZN(new_n405));
  INV_X1    g219(.A(G902), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n392), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n408), .B(KEYINPUT91), .Z(new_n410));
  AOI22_X1  g224(.A1(new_n365), .A2(new_n368), .B1(new_n389), .B2(new_n390), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n406), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n332), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n241), .A2(G122), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT14), .Z(new_n416));
  INV_X1    g230(.A(G122), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G116), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT94), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G107), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n337), .A3(new_n415), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n191), .A2(G128), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n196), .A2(G143), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(G134), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT95), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n421), .A2(new_n429), .A3(new_n422), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n419), .A2(new_n415), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G107), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n422), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n216), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(new_n425), .Z(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT9), .B(G234), .ZN(new_n439));
  INV_X1    g253(.A(G217), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(G953), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n431), .B2(new_n438), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n406), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G478), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n447), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G113), .B(G122), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(new_n334), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n270), .A2(G143), .A3(G214), .ZN(new_n453));
  AOI21_X1  g267(.A(G143), .B1(new_n270), .B2(G214), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n210), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT18), .ZN(new_n457));
  XNOR2_X1  g271(.A(G125), .B(G140), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(new_n189), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT92), .B1(new_n460), .B2(new_n210), .ZN(new_n461));
  OR3_X1    g275(.A1(new_n460), .A2(new_n210), .A3(KEYINPUT92), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n455), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(KEYINPUT16), .ZN(new_n465));
  OR3_X1    g279(.A1(new_n370), .A2(KEYINPUT16), .A3(G140), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(G146), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n455), .B(new_n210), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT17), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n452), .B(new_n464), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(G146), .A3(new_n466), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n458), .B(KEYINPUT19), .Z(new_n476));
  OAI211_X1 g290(.A(new_n471), .B(new_n475), .C1(G146), .C2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n452), .B1(new_n477), .B2(new_n464), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(G475), .A2(G902), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT93), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT20), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n477), .A2(new_n464), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n473), .B1(new_n484), .B2(new_n452), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n481), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n470), .A2(new_n472), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n452), .B1(new_n489), .B2(new_n464), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n406), .B1(new_n490), .B2(new_n474), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(G234), .A2(G237), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n494), .A2(G952), .A3(new_n386), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n494), .A2(G902), .A3(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT21), .B(G898), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n450), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n414), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT80), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n198), .A2(new_n354), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n195), .A2(new_n197), .A3(new_n343), .A4(new_n353), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n215), .A2(new_n278), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n504), .B2(KEYINPUT12), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT80), .B(new_n506), .C1(new_n507), .C2(new_n230), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(KEYINPUT12), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT79), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n280), .A2(new_n511), .A3(new_n344), .A4(new_n346), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n254), .A2(new_n258), .A3(new_n346), .ZN(new_n513));
  INV_X1    g327(.A(new_n344), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT79), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n503), .B(KEYINPUT10), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n230), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G140), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n386), .A2(G227), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n517), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n279), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n522), .A3(new_n518), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n527), .A3(G469), .ZN(new_n528));
  INV_X1    g342(.A(G469), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(new_n406), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n510), .A2(new_n518), .A3(new_n522), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT82), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n510), .A2(new_n518), .A3(new_n535), .A4(new_n522), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n526), .A2(new_n518), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT81), .B(G469), .Z(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n406), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT83), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n534), .A2(new_n536), .B1(new_n523), .B2(new_n538), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G902), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT83), .A3(new_n541), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n532), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G221), .ZN(new_n549));
  INV_X1    g363(.A(new_n439), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n406), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n500), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT23), .B1(new_n196), .B2(G119), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT77), .B1(new_n239), .B2(G128), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n553), .B(new_n554), .Z(new_n555));
  AND2_X1   g369(.A1(new_n555), .A2(G110), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  XNOR2_X1  g371(.A(G119), .B(G128), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OR3_X1    g373(.A1(new_n468), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n555), .A2(G110), .B1(new_n558), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n458), .A2(new_n189), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n475), .A3(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT22), .B(G137), .Z(new_n564));
  NAND3_X1  g378(.A1(new_n386), .A2(G221), .A3(G234), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n560), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n560), .B2(new_n563), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n440), .B1(G234), .B2(new_n406), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n406), .B1(new_n567), .B2(new_n568), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT25), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(new_n570), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n330), .A2(new_n552), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(G101), .ZN(G3));
  OAI21_X1  g394(.A(G472), .B1(new_n299), .B2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n302), .A2(new_n581), .A3(new_n308), .ZN(new_n582));
  INV_X1    g396(.A(new_n578), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n548), .A2(new_n551), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n408), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n411), .B2(new_n412), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n409), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n331), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n445), .A2(G478), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT33), .B1(new_n443), .B2(new_n444), .ZN(new_n592));
  INV_X1    g406(.A(new_n444), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n442), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n493), .B(new_n591), .C1(new_n596), .C2(new_n446), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n590), .A2(new_n498), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n586), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT96), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(KEYINPUT97), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT98), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n601), .B(new_n603), .ZN(G6));
  AOI21_X1  g418(.A(new_n332), .B1(new_n409), .B2(new_n588), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n450), .A2(new_n492), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n487), .A2(KEYINPUT99), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(new_n483), .Z(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n498), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n586), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G107), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  INV_X1    g428(.A(new_n582), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n577), .A2(new_n570), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n560), .A2(new_n563), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n571), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n552), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  INV_X1    g438(.A(G900), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n495), .B1(new_n496), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n616), .A2(new_n620), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n590), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n330), .A2(new_n585), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n330), .A2(KEYINPUT100), .A3(new_n630), .A4(new_n585), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G128), .ZN(G30));
  NAND2_X1  g450(.A1(new_n409), .A2(new_n413), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n409), .A2(new_n413), .A3(KEYINPUT38), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n483), .A2(new_n487), .B1(G475), .B2(new_n491), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n449), .B2(new_n448), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n629), .A2(new_n331), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n626), .B(KEYINPUT39), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n585), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n641), .B(new_n644), .C1(new_n646), .C2(KEYINPUT40), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n648));
  INV_X1    g462(.A(new_n319), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n649), .A2(new_n275), .B1(new_n294), .B2(new_n297), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT101), .B(G143), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G45));
  NOR2_X1   g470(.A1(new_n597), .A2(new_n626), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n605), .A2(new_n657), .A3(new_n621), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n330), .A2(new_n585), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n551), .ZN(new_n661));
  OAI21_X1  g475(.A(G469), .B1(new_n545), .B2(G902), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT83), .B1(new_n546), .B2(new_n541), .ZN(new_n663));
  INV_X1    g477(.A(new_n541), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n545), .A2(new_n543), .A3(G902), .A4(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n330), .A2(new_n578), .A3(new_n598), .A4(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NAND4_X1  g488(.A1(new_n330), .A2(new_n611), .A3(new_n578), .A4(new_n667), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NOR2_X1   g490(.A1(new_n666), .A2(new_n590), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n499), .A3(new_n621), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n330), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G119), .ZN(G21));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n275), .A2(new_n320), .B1(new_n289), .B2(new_n298), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(new_n301), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n320), .A2(new_n275), .ZN(new_n684));
  OAI211_X1 g498(.A(KEYINPUT103), .B(new_n300), .C1(new_n684), .C2(new_n306), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n578), .A3(new_n581), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n605), .A2(new_n610), .A3(new_n643), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n687), .A2(new_n688), .A3(new_n666), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n417), .ZN(G24));
  AND4_X1   g504(.A1(new_n581), .A2(new_n686), .A3(new_n621), .A4(new_n657), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n677), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  NAND3_X1  g507(.A1(new_n409), .A2(new_n413), .A3(new_n331), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n528), .A2(KEYINPUT104), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n528), .A2(KEYINPUT104), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n531), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n544), .B2(new_n547), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n551), .ZN(new_n701));
  INV_X1    g515(.A(new_n697), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n528), .A2(KEYINPUT104), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n530), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n663), .B2(new_n665), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT105), .B1(new_n705), .B2(new_n661), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n695), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n313), .B(KEYINPUT32), .ZN(new_n708));
  INV_X1    g522(.A(new_n329), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n578), .B(new_n657), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT42), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n700), .B1(new_n699), .B2(new_n551), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n705), .A2(KEYINPUT105), .A3(new_n661), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n694), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n597), .A2(KEYINPUT42), .A3(new_n626), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n330), .A3(new_n578), .A4(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  INV_X1    g532(.A(new_n628), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n330), .A3(new_n578), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  OAI211_X1 g535(.A(new_n591), .B(new_n642), .C1(new_n596), .C2(new_n446), .ZN(new_n722));
  NOR2_X1   g536(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n722), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n582), .A3(new_n621), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n524), .A2(new_n527), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n731), .B(G469), .C1(new_n734), .C2(G902), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n732), .A2(new_n733), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n531), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n544), .A2(new_n547), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n661), .A3(new_n645), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n727), .A2(KEYINPUT44), .A3(new_n582), .A4(new_n621), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n730), .A2(new_n742), .A3(new_n695), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  NAND2_X1  g559(.A1(new_n741), .A2(new_n661), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n741), .A2(KEYINPUT47), .A3(new_n661), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n330), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n694), .A2(new_n578), .A3(new_n597), .A4(new_n626), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT107), .B(G140), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G42));
  INV_X1    g569(.A(new_n652), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n740), .A2(new_n662), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT49), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n583), .A2(new_n551), .A3(new_n332), .A4(new_n722), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n756), .A2(new_n641), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n689), .B1(new_n678), .B2(new_n330), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n675), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n670), .B2(new_n671), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n414), .A2(new_n610), .ZN(new_n764));
  INV_X1    g578(.A(new_n597), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n584), .A2(new_n764), .A3(new_n585), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n579), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT108), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n579), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n606), .B1(new_n483), .B2(new_n487), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n584), .A2(new_n764), .A3(new_n585), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n622), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n768), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n448), .A2(new_n449), .A3(new_n492), .A4(new_n627), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT109), .B1(new_n608), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n621), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n608), .A2(new_n776), .A3(KEYINPUT109), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n694), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n330), .A2(new_n585), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n691), .B(new_n695), .C1(new_n706), .C2(new_n701), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n711), .A3(new_n716), .A4(new_n720), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n775), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n659), .A2(new_n692), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n633), .B2(new_n634), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n605), .A2(new_n643), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n788), .A2(new_n629), .A3(new_n627), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n652), .A2(new_n661), .A3(new_n705), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n786), .ZN(new_n792));
  AND4_X1   g606(.A1(KEYINPUT52), .A2(new_n635), .A3(new_n792), .A4(new_n790), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n763), .B(new_n785), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n773), .B1(new_n767), .B2(KEYINPUT108), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n720), .A2(new_n782), .A3(new_n781), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n717), .A3(new_n799), .A4(new_n770), .ZN(new_n800));
  INV_X1    g614(.A(new_n762), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n672), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n635), .A2(new_n792), .A3(new_n790), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n787), .A2(KEYINPUT52), .A3(new_n790), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n808), .A3(KEYINPUT53), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n796), .A2(new_n797), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n687), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n495), .A3(new_n727), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n331), .B1(new_n639), .B2(new_n640), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n667), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n815), .A3(KEYINPUT114), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n495), .A3(new_n727), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n814), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(KEYINPUT115), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n812), .A2(new_n815), .A3(KEYINPUT50), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n823), .A2(KEYINPUT115), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n816), .B2(new_n819), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n666), .A2(new_n694), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n578), .A3(new_n495), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n652), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n596), .A2(new_n446), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n493), .B1(new_n830), .B2(new_n591), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n495), .A3(new_n727), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n686), .A2(new_n581), .A3(new_n621), .ZN(new_n833));
  OR3_X1    g647(.A1(new_n832), .A2(KEYINPUT116), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n829), .A2(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(KEYINPUT117), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n826), .B2(new_n836), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n757), .A2(new_n551), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n750), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n818), .A2(new_n694), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT112), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n843), .B1(new_n750), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n840), .A2(new_n842), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n386), .A2(G952), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n852), .B1(new_n812), .B2(new_n677), .ZN(new_n853));
  INV_X1    g667(.A(new_n829), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n597), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n853), .B(KEYINPUT119), .C1(new_n854), .C2(new_n597), .ZN(new_n858));
  AND2_X1   g672(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n708), .A2(new_n709), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n832), .A2(new_n860), .A3(new_n583), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n844), .B(KEYINPUT113), .Z(new_n865));
  OAI21_X1  g679(.A(new_n848), .B1(new_n750), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n826), .A2(new_n836), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n837), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n851), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n796), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n803), .B2(new_n808), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT110), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n809), .A2(KEYINPUT111), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n803), .A2(new_n808), .A3(new_n875), .A4(KEYINPUT53), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n810), .B(new_n869), .C1(new_n877), .C2(KEYINPUT54), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n760), .B1(new_n878), .B2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n796), .A2(new_n809), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(G902), .A3(new_n410), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n369), .A2(new_n391), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n411), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n882), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n386), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n406), .B1(new_n796), .B2(new_n809), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(new_n587), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(new_n885), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n896), .ZN(G51));
  XNOR2_X1  g711(.A(new_n530), .B(KEYINPUT57), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n797), .B1(new_n796), .B2(new_n809), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n810), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n540), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(G469), .A3(new_n734), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n892), .B1(new_n901), .B2(new_n902), .ZN(G54));
  NAND2_X1  g717(.A1(KEYINPUT58), .A2(G475), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n894), .A2(new_n485), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n485), .B1(new_n894), .B2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n892), .ZN(G60));
  INV_X1    g722(.A(new_n592), .ZN(new_n909));
  INV_X1    g723(.A(new_n595), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT59), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n912), .B(new_n914), .C1(new_n810), .C2(new_n899), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n893), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n874), .A2(new_n876), .ZN(new_n917));
  AOI211_X1 g731(.A(new_n870), .B(KEYINPUT53), .C1(new_n803), .C2(new_n808), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT110), .B1(new_n794), .B2(new_n795), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n797), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n921), .B2(new_n810), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n916), .B1(new_n922), .B2(new_n911), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  NAND2_X1  g739(.A1(new_n881), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n569), .B(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n881), .A2(new_n619), .A3(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n893), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(G66));
  NAND3_X1  g748(.A1(new_n763), .A2(new_n770), .A3(new_n798), .ZN(new_n935));
  NAND2_X1  g749(.A1(G224), .A2(G953), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n935), .A2(G953), .B1(new_n497), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n365), .B(new_n368), .C1(G898), .C2(new_n386), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n937), .B(new_n938), .Z(G69));
  NOR2_X1   g753(.A1(new_n277), .A2(new_n282), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n476), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(G900), .B2(G953), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n860), .A2(new_n583), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n788), .A3(new_n742), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n720), .A2(new_n753), .A3(new_n744), .A4(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n717), .A3(new_n787), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n945), .A2(new_n948), .A3(new_n717), .A4(new_n787), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n942), .B1(new_n950), .B2(G953), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n695), .B1(new_n771), .B2(new_n765), .ZN(new_n952));
  OR4_X1    g766(.A1(new_n751), .A2(new_n583), .A3(new_n646), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n744), .A3(new_n753), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n654), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n957), .B(new_n787), .C1(new_n958), .C2(KEYINPUT62), .ZN(new_n959));
  INV_X1    g773(.A(new_n787), .ZN(new_n960));
  OAI211_X1 g774(.A(KEYINPUT123), .B(new_n955), .C1(new_n960), .C2(new_n654), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n954), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n941), .B1(new_n962), .B2(G953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n386), .B1(G227), .B2(G900), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n951), .A2(new_n963), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n965), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(G72));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n950), .B2(new_n935), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n892), .B1(new_n976), .B2(new_n326), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  INV_X1    g792(.A(new_n935), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n978), .B1(new_n962), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n325), .A2(new_n274), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n325), .A2(new_n275), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n294), .A2(new_n297), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n877), .A2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n877), .A2(KEYINPUT127), .A3(new_n985), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(G57));
endmodule


