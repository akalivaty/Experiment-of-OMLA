//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  INV_X1    g002(.A(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT75), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT74), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n212), .ZN(new_n214));
  AND4_X1   g013(.A1(new_n207), .A2(new_n213), .A3(new_n210), .A4(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n206), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n210), .A3(new_n214), .ZN(new_n217));
  INV_X1    g016(.A(new_n207), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n209), .A2(new_n207), .A3(new_n210), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT77), .B(G162gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n233), .A2(new_n235), .B1(new_n223), .B2(new_n224), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n227), .B(new_n228), .C1(new_n231), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n216), .A2(new_n221), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G228gat), .ZN(new_n243));
  INV_X1    g042(.A(G233gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n227), .B1(new_n231), .B2(new_n236), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n219), .B2(new_n220), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n247), .B2(KEYINPUT3), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n216), .A2(KEYINPUT80), .A3(new_n239), .A4(new_n221), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n245), .A3(new_n248), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n219), .A2(new_n220), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n238), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(KEYINPUT78), .ZN(new_n254));
  INV_X1    g053(.A(G162gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT77), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT77), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G162gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(G155gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT2), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n234), .A2(G141gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n232), .A2(G148gat), .ZN(new_n262));
  INV_X1    g061(.A(G155gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n255), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n261), .A2(new_n262), .B1(new_n264), .B2(new_n222), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n229), .B1(new_n233), .B2(new_n235), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n260), .A2(new_n265), .B1(new_n266), .B2(new_n225), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n253), .A2(new_n228), .B1(new_n254), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n252), .B1(new_n237), .B2(new_n238), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n270), .A2(new_n271), .B1(new_n243), .B2(new_n244), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n250), .A2(new_n251), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n251), .B1(new_n250), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G22gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n250), .A2(new_n272), .A3(new_n251), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n205), .A2(KEYINPUT81), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(KEYINPUT81), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n275), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT35), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(G127gat), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT69), .B(G134gat), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n289), .B2(G134gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n287), .A3(G127gat), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  INV_X1    g097(.A(G113gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G120gat), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G113gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT70), .B1(new_n299), .B2(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n301), .A3(G113gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n302), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT1), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n287), .A2(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n289), .A2(G134gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n304), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT27), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G183gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT27), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(G183gat), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT66), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT28), .A3(new_n319), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(G169gat), .ZN(new_n334));
  INV_X1    g133(.A(G176gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n334), .A3(new_n335), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n342), .A2(new_n343), .B1(G169gat), .B2(G176gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n332), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n346), .B(new_n347), .C1(G183gat), .C2(G190gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT25), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(new_n324), .A3(new_n319), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n346), .A3(new_n347), .A4(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n317), .A2(new_n340), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G227gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n244), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n297), .A2(new_n303), .B1(new_n309), .B2(new_n315), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n344), .A2(new_n348), .A3(KEYINPUT25), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n344), .B2(new_n353), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n338), .B1(new_n328), .B2(new_n330), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n357), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT32), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT72), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(G71gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(G99gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n374), .A3(KEYINPUT32), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n368), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n366), .B(KEYINPUT32), .C1(new_n372), .C2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n365), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n358), .B2(new_n244), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n380), .A2(KEYINPUT34), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(KEYINPUT34), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n376), .A2(new_n382), .A3(new_n377), .A4(new_n381), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n283), .A2(new_n284), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  INV_X1    g187(.A(G64gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G92gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n340), .A2(new_n356), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n340), .B2(new_n356), .ZN(new_n398));
  INV_X1    g197(.A(new_n252), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n216), .A2(new_n221), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n238), .B1(new_n363), .B2(new_n364), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(new_n398), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n392), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n363), .A2(new_n364), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n393), .B1(new_n407), .B2(KEYINPUT29), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(new_n404), .A3(new_n252), .ZN(new_n409));
  INV_X1    g208(.A(new_n392), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n393), .B2(new_n402), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n401), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n412), .A3(KEYINPUT30), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n400), .A2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT30), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n410), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n360), .A2(KEYINPUT4), .A3(new_n254), .A4(new_n269), .ZN(new_n418));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT4), .ZN(new_n420));
  INV_X1    g219(.A(new_n237), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n260), .A2(new_n265), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n228), .B1(new_n422), .B2(new_n227), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n420), .B1(new_n424), .B2(new_n317), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n304), .A2(new_n267), .A3(new_n316), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n418), .B(new_n419), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n317), .A2(new_n246), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n426), .ZN(new_n430));
  INV_X1    g229(.A(new_n419), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(KEYINPUT5), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n424), .A2(new_n317), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(KEYINPUT4), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n360), .A2(new_n420), .A3(new_n254), .A4(new_n269), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT79), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT79), .B1(new_n436), .B2(new_n437), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n434), .B(new_n435), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G1gat), .B(G29gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT0), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G57gat), .ZN(new_n444));
  INV_X1    g243(.A(G85gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n440), .A3(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n417), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n387), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n384), .A2(new_n458), .A3(new_n385), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n378), .A2(KEYINPUT73), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n282), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n457), .B(new_n284), .C1(new_n461), .C2(new_n453), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n459), .A2(new_n460), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n453), .A3(new_n283), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT82), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n456), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n459), .B2(new_n460), .ZN(new_n469));
  OR2_X1    g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n414), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n400), .B2(new_n405), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n392), .A3(new_n473), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n474), .A2(KEYINPUT38), .B1(new_n414), .B2(new_n410), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n411), .A2(new_n401), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n252), .B1(new_n408), .B2(new_n404), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT37), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n478), .A3(new_n479), .A4(new_n392), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(new_n452), .A3(new_n451), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n436), .A2(new_n437), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT79), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n484), .A2(new_n485), .B1(new_n424), .B2(new_n317), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(new_n419), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n447), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n429), .A2(new_n419), .A3(new_n426), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT39), .B(new_n490), .C1(new_n486), .C2(new_n419), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n448), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n417), .B1(new_n492), .B2(new_n493), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n283), .B(new_n481), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n470), .B(new_n497), .C1(new_n453), .C2(new_n283), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n466), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT84), .ZN(new_n503));
  XOR2_X1   g302(.A(G113gat), .B(G141gat), .Z(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G169gat), .B(G197gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT12), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT16), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n511), .B(new_n512), .C1(new_n510), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g312(.A1(KEYINPUT87), .A2(G8gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT14), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n204), .A2(G43gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(KEYINPUT85), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n520), .B(new_n523), .C1(new_n524), .C2(new_n519), .ZN(new_n525));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n519), .A2(new_n524), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n519), .B2(new_n518), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n525), .B(new_n526), .C1(new_n529), .C2(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT86), .A2(KEYINPUT17), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n527), .A2(new_n530), .A3(new_n533), .A4(new_n534), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n515), .A2(new_n531), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n515), .B(new_n531), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n540), .B(KEYINPUT13), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n508), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n538), .A2(new_n539), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(KEYINPUT18), .ZN(new_n552));
  AND4_X1   g351(.A1(new_n508), .A2(new_n551), .A3(new_n547), .A4(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n501), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n544), .A2(new_n508), .A3(new_n547), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n547), .A3(new_n552), .ZN(new_n556));
  INV_X1    g355(.A(new_n508), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n558), .A3(KEYINPUT88), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n500), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G57gat), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n567), .A2(new_n389), .A3(KEYINPUT90), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n389), .B1(new_n567), .B2(KEYINPUT90), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n563), .B(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT91), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n515), .B1(new_n578), .B2(KEYINPUT21), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G127gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  XNOR2_X1  g383(.A(G155gat), .B(G183gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n583), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  INV_X1    g387(.A(G211gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n590), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n445), .B2(new_n391), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n596), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n531), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n536), .A2(new_n537), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n602), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT93), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n606), .A2(new_n608), .ZN(new_n610));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT94), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n609), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n615), .B1(new_n609), .B2(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n244), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621));
  INV_X1    g420(.A(new_n576), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT95), .B1(new_n598), .B2(new_n600), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n598), .A2(KEYINPUT95), .A3(new_n600), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n596), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n594), .B(KEYINPUT92), .ZN(new_n629));
  INV_X1    g428(.A(new_n625), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(new_n623), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n631), .A2(KEYINPUT96), .B1(new_n629), .B2(new_n601), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n621), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(new_n601), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n626), .B2(new_n627), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n576), .B1(new_n631), .B2(KEYINPUT96), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(KEYINPUT97), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n602), .A2(new_n622), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n633), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n578), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT98), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n578), .A2(new_n643), .A3(KEYINPUT10), .A4(new_n602), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n620), .B1(new_n640), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n633), .A2(new_n639), .A3(new_n637), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n620), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n335), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(G204gat), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n593), .A2(new_n618), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n562), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT99), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n451), .A2(new_n452), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n662), .ZN(new_n667));
  INV_X1    g466(.A(new_n417), .ZN(new_n668));
  OAI21_X1  g467(.A(G8gat), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OR2_X1    g469(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n662), .A2(new_n417), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(new_n670), .ZN(new_n676));
  OAI221_X1 g475(.A(new_n669), .B1(new_n670), .B2(new_n673), .C1(new_n675), .C2(new_n676), .ZN(G1325gat));
  AOI21_X1  g476(.A(G15gat), .B1(new_n662), .B2(new_n386), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n667), .A2(new_n470), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n662), .A2(new_n282), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  INV_X1    g483(.A(new_n618), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n499), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n457), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n464), .A2(KEYINPUT82), .A3(KEYINPUT35), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n455), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n453), .B2(new_n283), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n454), .A2(KEYINPUT101), .A3(new_n282), .ZN(new_n693));
  AND4_X1   g492(.A1(new_n470), .A2(new_n497), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n684), .B(new_n685), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n470), .A2(new_n497), .A3(new_n692), .A4(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n618), .B1(new_n466), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(KEYINPUT102), .A3(new_n684), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n686), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n593), .A2(new_n657), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n548), .A2(new_n553), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n701), .A2(KEYINPUT103), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  INV_X1    g506(.A(new_n686), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n466), .A2(new_n698), .ZN(new_n709));
  AND4_X1   g508(.A1(KEYINPUT102), .A2(new_n709), .A3(new_n684), .A4(new_n685), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT102), .B1(new_n699), .B2(new_n684), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n705), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n663), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n562), .A2(new_n685), .A3(new_n702), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n516), .A3(new_n664), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1328gat));
  OAI21_X1  g519(.A(G36gat), .B1(new_n715), .B2(new_n668), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT46), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n717), .A2(new_n517), .A3(new_n417), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(KEYINPUT46), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(new_n470), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n706), .B2(new_n714), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT103), .B1(new_n701), .B2(new_n705), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n712), .A2(new_n707), .A3(new_n713), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n470), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n735), .A3(new_n386), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n731), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n712), .A2(new_n713), .ZN(new_n741));
  OAI21_X1  g540(.A(G43gat), .B1(new_n741), .B2(new_n470), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n737), .A3(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1330gat));
  OAI21_X1  g543(.A(G50gat), .B1(new_n741), .B2(new_n283), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n717), .A2(new_n204), .A3(new_n282), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT48), .ZN(new_n747));
  OAI21_X1  g546(.A(G50gat), .B1(new_n715), .B2(new_n283), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n746), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g549(.A(new_n704), .B1(new_n466), .B2(new_n698), .ZN(new_n751));
  INV_X1    g550(.A(new_n593), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n685), .A3(new_n658), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n663), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n567), .ZN(G1332gat));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n668), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754), .B2(new_n470), .ZN(new_n762));
  INV_X1    g561(.A(new_n386), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(G71gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n754), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n754), .A2(new_n283), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n703), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n701), .A2(new_n658), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n664), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n699), .A2(new_n703), .A3(new_n752), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT106), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n664), .A2(new_n445), .A3(new_n657), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT107), .Z(new_n780));
  OAI22_X1  g579(.A1(new_n771), .A2(new_n445), .B1(new_n778), .B2(new_n780), .ZN(G1336gat));
  NAND2_X1  g580(.A1(new_n770), .A2(new_n417), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G92gat), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n658), .A2(G92gat), .A3(new_n668), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n783), .B(new_n784), .C1(new_n778), .C2(new_n786), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n782), .A2(KEYINPUT108), .A3(G92gat), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT108), .B1(new_n782), .B2(G92gat), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n785), .B(KEYINPUT109), .Z(new_n790));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n792), .B2(new_n784), .ZN(G1337gat));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n774), .A2(new_n777), .A3(new_n795), .A4(new_n657), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n763), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n770), .A2(new_n728), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI221_X1 g599(.A(KEYINPUT110), .B1(new_n798), .B2(new_n795), .C1(new_n796), .C2(new_n763), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1338gat));
  NAND2_X1  g601(.A1(new_n770), .A2(new_n282), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n658), .A2(G106gat), .A3(new_n283), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n804), .B(new_n805), .C1(new_n778), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n773), .A2(new_n807), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n803), .B2(G106gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n805), .ZN(G1339gat));
  NOR2_X1   g610(.A1(new_n663), .A2(new_n417), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n655), .B1(new_n646), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n640), .A2(new_n645), .A3(new_n620), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n646), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n817), .B2(KEYINPUT54), .ZN(new_n818));
  NOR4_X1   g617(.A1(new_n816), .A2(new_n646), .A3(KEYINPUT112), .A4(new_n813), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n814), .B(KEYINPUT55), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n704), .A3(new_n656), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n549), .A2(new_n540), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n826), .B(new_n827), .C1(new_n545), .C2(new_n546), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n553), .B1(new_n828), .B2(new_n507), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n657), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n685), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n822), .A2(new_n656), .A3(new_n823), .A4(new_n829), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n618), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n752), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT111), .B1(new_n660), .B2(new_n703), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n659), .A2(new_n836), .A3(new_n704), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n282), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n386), .B(new_n812), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843), .B2(new_n561), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n663), .B1(new_n834), .B2(new_n838), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(new_n668), .A3(new_n461), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n299), .A3(new_n704), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n843), .B2(new_n658), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n301), .A3(new_n657), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  INV_X1    g650(.A(new_n843), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n286), .A3(new_n593), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n286), .B1(new_n846), .B2(new_n593), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1342gat));
  NAND3_X1  g657(.A1(new_n846), .A2(new_n287), .A3(new_n685), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n859), .B(KEYINPUT56), .Z(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n843), .B2(new_n618), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n860), .A2(KEYINPUT116), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1343gat));
  NAND2_X1  g665(.A1(new_n834), .A2(new_n838), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n664), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n561), .A2(G141gat), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n728), .A2(new_n283), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n668), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n870), .A2(new_n871), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT119), .B1(new_n867), .B2(new_n664), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n869), .B(new_n663), .C1(new_n834), .C2(new_n838), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n871), .A4(new_n874), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n470), .A2(new_n812), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT117), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n822), .A2(new_n560), .A3(new_n656), .A4(new_n823), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n685), .B1(new_n887), .B2(new_n830), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n752), .B1(new_n888), .B2(new_n833), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT118), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n891), .B(new_n752), .C1(new_n888), .C2(new_n833), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n838), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n283), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n867), .A2(new_n282), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n894), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n886), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n232), .B1(new_n899), .B2(new_n704), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT58), .B1(new_n883), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n879), .A2(new_n880), .A3(new_n873), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT58), .B1(new_n902), .B2(new_n871), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n899), .A2(new_n560), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n232), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT121), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n902), .A2(new_n234), .A3(new_n657), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT57), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n889), .B1(new_n560), .B2(new_n659), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n894), .A3(new_n282), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n657), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n885), .B(KEYINPUT122), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n234), .C1(new_n899), .C2(new_n657), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n911), .B1(new_n919), .B2(new_n920), .ZN(G1345gat));
  AOI21_X1  g720(.A(G155gat), .B1(new_n902), .B2(new_n593), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n752), .A2(new_n263), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n899), .B2(new_n923), .ZN(G1346gat));
  INV_X1    g723(.A(new_n230), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n925), .A3(new_n685), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n685), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(new_n925), .ZN(G1347gat));
  OR2_X1    g728(.A1(new_n841), .A2(new_n842), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n664), .A2(new_n668), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n386), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT125), .Z(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n560), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G169gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n867), .A2(new_n663), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT124), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(new_n417), .A3(new_n461), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n704), .A2(new_n334), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  NAND4_X1  g739(.A1(new_n930), .A2(G176gat), .A3(new_n657), .A4(new_n933), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n938), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n657), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n944), .B2(new_n335), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n329), .A3(new_n593), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n593), .A3(new_n933), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G183gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n943), .A2(new_n319), .A3(new_n685), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n930), .A2(new_n685), .A3(new_n933), .ZN(new_n955));
  XOR2_X1   g754(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n955), .A2(G190gat), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n955), .B2(G190gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NAND4_X1  g759(.A1(new_n913), .A2(new_n470), .A3(new_n915), .A4(new_n931), .ZN(new_n961));
  OAI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n561), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n937), .A2(new_n872), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n417), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n703), .A2(G197gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  XNOR2_X1  g765(.A(KEYINPUT127), .B(G204gat), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n963), .A2(new_n417), .A3(new_n657), .A4(new_n968), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n470), .A2(new_n931), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n916), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n969), .A2(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(G1353gat));
  INV_X1    g773(.A(new_n964), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n589), .A3(new_n593), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n961), .A2(new_n752), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n961), .A2(new_n981), .A3(new_n618), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n975), .A2(new_n685), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n983), .B2(new_n981), .ZN(G1355gat));
endmodule


