

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727;

  XNOR2_X1 U368 ( .A(n711), .B(G146), .ZN(n507) );
  NOR2_X2 U369 ( .A1(G902), .A2(n679), .ZN(n510) );
  NOR2_X1 U370 ( .A1(n727), .A2(n722), .ZN(n542) );
  INV_X1 U371 ( .A(G953), .ZN(n714) );
  NOR2_X2 U372 ( .A1(n394), .A2(n591), .ZN(n576) );
  XNOR2_X2 U373 ( .A(n417), .B(n471), .ZN(n569) );
  NAND2_X1 U374 ( .A1(n726), .A2(n612), .ZN(n579) );
  AND2_X1 U375 ( .A1(n583), .A2(n353), .ZN(n408) );
  XNOR2_X1 U376 ( .A(n363), .B(KEYINPUT112), .ZN(n725) );
  XNOR2_X1 U377 ( .A(n392), .B(KEYINPUT22), .ZN(n431) );
  XNOR2_X1 U378 ( .A(n508), .B(G469), .ZN(n509) );
  INV_X1 U379 ( .A(n551), .ZN(n346) );
  XNOR2_X1 U380 ( .A(n393), .B(n355), .ZN(n558) );
  XNOR2_X1 U381 ( .A(n374), .B(n354), .ZN(n711) );
  OR2_X1 U382 ( .A1(G902), .A2(G237), .ZN(n525) );
  XNOR2_X1 U383 ( .A(n542), .B(KEYINPUT46), .ZN(n366) );
  XNOR2_X1 U384 ( .A(n441), .B(n473), .ZN(n442) );
  XNOR2_X1 U385 ( .A(G110), .B(G104), .ZN(n500) );
  XNOR2_X1 U386 ( .A(n524), .B(n707), .ZN(n671) );
  XNOR2_X1 U387 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U388 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U389 ( .A(n374), .B(n429), .ZN(n523) );
  NOR2_X1 U390 ( .A1(n380), .A2(n378), .ZN(n377) );
  NAND2_X1 U391 ( .A1(n379), .A2(n350), .ZN(n378) );
  NOR2_X1 U392 ( .A1(n663), .A2(n381), .ZN(n380) );
  XNOR2_X1 U393 ( .A(n571), .B(KEYINPUT106), .ZN(n391) );
  NOR2_X1 U394 ( .A1(G953), .A2(G237), .ZN(n465) );
  NAND2_X1 U395 ( .A1(n371), .A2(n369), .ZN(n561) );
  AND2_X1 U396 ( .A1(n549), .A2(n351), .ZN(n371) );
  INV_X1 U397 ( .A(KEYINPUT107), .ZN(n389) );
  XNOR2_X1 U398 ( .A(G113), .B(KEYINPUT3), .ZN(n460) );
  XNOR2_X1 U399 ( .A(G119), .B(G116), .ZN(n462) );
  INV_X1 U400 ( .A(KEYINPUT44), .ZN(n580) );
  INV_X1 U401 ( .A(KEYINPUT1), .ZN(n511) );
  NAND2_X1 U402 ( .A1(n424), .A2(n423), .ZN(n636) );
  INV_X1 U403 ( .A(n564), .ZN(n423) );
  NAND2_X1 U404 ( .A1(n352), .A2(n566), .ZN(n427) );
  OR2_X1 U405 ( .A1(n597), .A2(G902), .ZN(n417) );
  XOR2_X1 U406 ( .A(G137), .B(G140), .Z(n501) );
  INV_X1 U407 ( .A(G101), .ZN(n502) );
  AND2_X1 U408 ( .A1(n725), .A2(n406), .ZN(n362) );
  XNOR2_X1 U409 ( .A(n420), .B(n419), .ZN(n534) );
  INV_X1 U410 ( .A(KEYINPUT39), .ZN(n419) );
  INV_X1 U411 ( .A(KEYINPUT19), .ZN(n428) );
  AND2_X1 U412 ( .A1(n585), .A2(n532), .ZN(n533) );
  INV_X1 U413 ( .A(n531), .ZN(n532) );
  XNOR2_X1 U414 ( .A(n372), .B(n457), .ZN(n555) );
  NOR2_X1 U415 ( .A1(n691), .A2(G902), .ZN(n372) );
  XNOR2_X1 U416 ( .A(n444), .B(n399), .ZN(n539) );
  XNOR2_X1 U417 ( .A(n445), .B(G475), .ZN(n399) );
  XNOR2_X1 U418 ( .A(n487), .B(n425), .ZN(n632) );
  XNOR2_X1 U419 ( .A(n486), .B(n426), .ZN(n425) );
  INV_X1 U420 ( .A(KEYINPUT25), .ZN(n426) );
  XNOR2_X1 U421 ( .A(n569), .B(n472), .ZN(n591) );
  INV_X1 U422 ( .A(KEYINPUT6), .ZN(n472) );
  XNOR2_X1 U423 ( .A(n516), .B(n405), .ZN(n707) );
  XNOR2_X1 U424 ( .A(n515), .B(n517), .ZN(n405) );
  NAND2_X1 U425 ( .A1(n370), .A2(n619), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n547), .B(KEYINPUT78), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n422), .B(G146), .ZN(n519) );
  INV_X1 U428 ( .A(G125), .ZN(n422) );
  AND2_X1 U429 ( .A1(n622), .A2(n625), .ZN(n651) );
  XOR2_X1 U430 ( .A(G131), .B(G122), .Z(n440) );
  XNOR2_X1 U431 ( .A(G113), .B(G104), .ZN(n439) );
  XNOR2_X1 U432 ( .A(G140), .B(G143), .ZN(n435) );
  XOR2_X1 U433 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n436) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n434) );
  XNOR2_X1 U435 ( .A(n519), .B(n421), .ZN(n473) );
  INV_X1 U436 ( .A(KEYINPUT10), .ZN(n421) );
  INV_X1 U437 ( .A(KEYINPUT4), .ZN(n459) );
  XNOR2_X1 U438 ( .A(n518), .B(n430), .ZN(n429) );
  INV_X1 U439 ( .A(KEYINPUT18), .ZN(n430) );
  INV_X1 U440 ( .A(n630), .ZN(n406) );
  AND2_X1 U441 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n463), .B(n464), .ZN(n516) );
  XNOR2_X1 U443 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U444 ( .A(KEYINPUT74), .ZN(n461) );
  XNOR2_X1 U445 ( .A(G122), .B(G134), .ZN(n447) );
  XNOR2_X1 U446 ( .A(n373), .B(KEYINPUT9), .ZN(n448) );
  INV_X1 U447 ( .A(KEYINPUT7), .ZN(n373) );
  XNOR2_X1 U448 ( .A(G116), .B(G107), .ZN(n450) );
  XNOR2_X1 U449 ( .A(n454), .B(n396), .ZN(n480) );
  XNOR2_X1 U450 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n396) );
  XOR2_X1 U451 ( .A(G902), .B(KEYINPUT15), .Z(n484) );
  XNOR2_X1 U452 ( .A(n540), .B(KEYINPUT41), .ZN(n664) );
  NAND2_X1 U453 ( .A1(n348), .A2(n640), .ZN(n644) );
  XNOR2_X1 U454 ( .A(n416), .B(n357), .ZN(n432) );
  OR2_X1 U455 ( .A1(n569), .A2(n529), .ZN(n416) );
  NOR2_X1 U456 ( .A1(n530), .A2(n636), .ZN(n585) );
  INV_X1 U457 ( .A(KEYINPUT89), .ZN(n567) );
  XNOR2_X1 U458 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U459 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U460 ( .A(n507), .B(n506), .ZN(n679) );
  XNOR2_X1 U461 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U462 ( .A(n673), .B(n672), .ZN(n674) );
  INV_X1 U463 ( .A(n693), .ZN(n698) );
  NAND2_X1 U464 ( .A1(n528), .A2(n551), .ZN(n363) );
  NAND2_X1 U465 ( .A1(n412), .A2(n410), .ZN(n727) );
  AND2_X1 U466 ( .A1(n413), .A2(n414), .ZN(n412) );
  NAND2_X1 U467 ( .A1(n411), .A2(n347), .ZN(n410) );
  NOR2_X1 U468 ( .A1(n550), .A2(n551), .ZN(n552) );
  INV_X1 U469 ( .A(KEYINPUT35), .ZN(n383) );
  NAND2_X1 U470 ( .A1(n391), .A2(n591), .ZN(n404) );
  NOR2_X1 U471 ( .A1(n640), .A2(n424), .ZN(n401) );
  INV_X1 U472 ( .A(n622), .ZN(n618) );
  AND2_X1 U473 ( .A1(n618), .A2(KEYINPUT40), .ZN(n347) );
  NOR2_X1 U474 ( .A1(n635), .A2(n636), .ZN(n348) );
  XNOR2_X1 U475 ( .A(n551), .B(KEYINPUT38), .ZN(n349) );
  INV_X1 U476 ( .A(n632), .ZN(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT80), .B(n578), .Z(n350) );
  OR2_X1 U478 ( .A1(KEYINPUT82), .A2(n548), .ZN(n351) );
  AND2_X1 U479 ( .A1(n631), .A2(n494), .ZN(n352) );
  AND2_X1 U480 ( .A1(n593), .A2(n604), .ZN(n353) );
  XOR2_X1 U481 ( .A(G131), .B(G134), .Z(n354) );
  XOR2_X1 U482 ( .A(n527), .B(n526), .Z(n355) );
  NOR2_X1 U483 ( .A1(n375), .A2(n640), .ZN(n356) );
  OR2_X1 U484 ( .A1(n539), .A2(n555), .ZN(n622) );
  XNOR2_X1 U485 ( .A(KEYINPUT113), .B(KEYINPUT30), .ZN(n357) );
  XOR2_X1 U486 ( .A(n577), .B(KEYINPUT81), .Z(n358) );
  XOR2_X1 U487 ( .A(n567), .B(KEYINPUT0), .Z(n359) );
  XOR2_X1 U488 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n360) );
  XNOR2_X1 U489 ( .A(n563), .B(KEYINPUT70), .ZN(n361) );
  XNOR2_X1 U490 ( .A(n365), .B(n361), .ZN(n364) );
  NAND2_X1 U491 ( .A1(n364), .A2(n362), .ZN(n713) );
  NAND2_X1 U492 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U493 ( .A(n562), .B(n368), .ZN(n367) );
  INV_X1 U494 ( .A(KEYINPUT71), .ZN(n368) );
  XNOR2_X2 U495 ( .A(n458), .B(n459), .ZN(n374) );
  OR2_X2 U496 ( .A1(n375), .A2(n568), .ZN(n392) );
  OR2_X1 U497 ( .A1(n375), .A2(n358), .ZN(n381) );
  NAND2_X1 U498 ( .A1(n375), .A2(n358), .ZN(n379) );
  NOR2_X1 U499 ( .A1(n375), .A2(n644), .ZN(n584) );
  XNOR2_X2 U500 ( .A(n400), .B(n359), .ZN(n375) );
  NAND2_X1 U501 ( .A1(n377), .A2(n376), .ZN(n382) );
  NAND2_X1 U502 ( .A1(n663), .A2(n358), .ZN(n376) );
  XNOR2_X2 U503 ( .A(n382), .B(n383), .ZN(n724) );
  NAND2_X1 U504 ( .A1(n385), .A2(n570), .ZN(n384) );
  NAND2_X1 U505 ( .A1(n386), .A2(n384), .ZN(n394) );
  NOR2_X1 U506 ( .A1(n636), .A2(n389), .ZN(n385) );
  NAND2_X1 U507 ( .A1(n636), .A2(n389), .ZN(n387) );
  NAND2_X1 U508 ( .A1(n635), .A2(n389), .ZN(n388) );
  XNOR2_X1 U509 ( .A(n498), .B(KEYINPUT109), .ZN(n499) );
  BUF_X1 U510 ( .A(n663), .Z(n390) );
  NAND2_X1 U511 ( .A1(n402), .A2(n401), .ZN(n612) );
  NAND2_X1 U512 ( .A1(n671), .A2(n595), .ZN(n393) );
  XNOR2_X1 U513 ( .A(n407), .B(n360), .ZN(n703) );
  NAND2_X1 U514 ( .A1(n581), .A2(n582), .ZN(n409) );
  NOR2_X1 U515 ( .A1(n695), .A2(G902), .ZN(n487) );
  XNOR2_X1 U516 ( .A(n483), .B(n395), .ZN(n695) );
  INV_X1 U517 ( .A(n710), .ZN(n395) );
  XNOR2_X1 U518 ( .A(n397), .B(KEYINPUT123), .ZN(G66) );
  NAND2_X1 U519 ( .A1(n699), .A2(n698), .ZN(n397) );
  NAND2_X1 U520 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U521 ( .A(n398), .B(n677), .ZN(G51) );
  NAND2_X1 U522 ( .A1(n676), .A2(n698), .ZN(n398) );
  NOR2_X2 U523 ( .A1(n565), .A2(n427), .ZN(n400) );
  XNOR2_X2 U524 ( .A(n543), .B(n428), .ZN(n565) );
  INV_X1 U525 ( .A(n590), .ZN(n402) );
  OR2_X1 U526 ( .A1(n431), .A2(n570), .ZN(n590) );
  XNOR2_X2 U527 ( .A(n403), .B(n572), .ZN(n726) );
  OR2_X2 U528 ( .A1(n431), .A2(n404), .ZN(n403) );
  NOR2_X1 U529 ( .A1(n703), .A2(n713), .ZN(n594) );
  XNOR2_X2 U530 ( .A(n446), .B(G143), .ZN(n458) );
  INV_X1 U531 ( .A(n534), .ZN(n411) );
  NAND2_X1 U532 ( .A1(n534), .A2(n415), .ZN(n413) );
  NAND2_X1 U533 ( .A1(n622), .A2(n415), .ZN(n414) );
  INV_X1 U534 ( .A(KEYINPUT40), .ZN(n415) );
  NAND2_X1 U535 ( .A1(n533), .A2(n432), .ZN(n556) );
  NAND2_X1 U536 ( .A1(n418), .A2(n533), .ZN(n420) );
  AND2_X1 U537 ( .A1(n432), .A2(n349), .ZN(n418) );
  INV_X1 U538 ( .A(KEYINPUT48), .ZN(n563) );
  INV_X1 U539 ( .A(KEYINPUT94), .ZN(n520) );
  XNOR2_X1 U540 ( .A(n467), .B(G137), .ZN(n468) );
  INV_X1 U541 ( .A(KEYINPUT104), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n574), .B(KEYINPUT108), .ZN(n575) );
  XNOR2_X1 U543 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U544 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U545 ( .A(n507), .B(n470), .ZN(n597) );
  XNOR2_X1 U546 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U547 ( .A(KEYINPUT105), .B(G478), .ZN(n457) );
  INV_X1 U548 ( .A(n695), .ZN(n696) );
  XOR2_X1 U549 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n514) );
  XNOR2_X1 U550 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n445) );
  NAND2_X1 U551 ( .A1(n465), .A2(G214), .ZN(n433) );
  XNOR2_X1 U552 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U553 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U554 ( .A(n438), .B(n437), .Z(n443) );
  XNOR2_X1 U555 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U556 ( .A(n443), .B(n442), .ZN(n684) );
  NOR2_X1 U557 ( .A1(G902), .A2(n684), .ZN(n444) );
  XNOR2_X2 U558 ( .A(G128), .B(KEYINPUT65), .ZN(n446) );
  XNOR2_X1 U559 ( .A(n448), .B(n447), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U561 ( .A(n458), .B(n453), .Z(n456) );
  NAND2_X1 U562 ( .A1(n714), .A2(G234), .ZN(n454) );
  NAND2_X1 U563 ( .A1(G217), .A2(n480), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n456), .B(n455), .ZN(n691) );
  XNOR2_X1 U565 ( .A(n460), .B(G101), .ZN(n464) );
  NAND2_X1 U566 ( .A1(n465), .A2(G210), .ZN(n466) );
  XNOR2_X1 U567 ( .A(n516), .B(n466), .ZN(n469) );
  XOR2_X1 U568 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n467) );
  XNOR2_X1 U569 ( .A(KEYINPUT77), .B(G472), .ZN(n471) );
  XOR2_X1 U570 ( .A(n501), .B(n473), .Z(n710) );
  XOR2_X1 U571 ( .A(KEYINPUT96), .B(G128), .Z(n475) );
  XNOR2_X1 U572 ( .A(G119), .B(G110), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n479) );
  XOR2_X1 U574 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n477) );
  XNOR2_X1 U575 ( .A(KEYINPUT79), .B(KEYINPUT85), .ZN(n476) );
  XNOR2_X1 U576 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U577 ( .A(n479), .B(n478), .Z(n482) );
  NAND2_X1 U578 ( .A1(G221), .A2(n480), .ZN(n481) );
  XNOR2_X1 U579 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U580 ( .A(KEYINPUT93), .B(n484), .ZN(n595) );
  NAND2_X1 U581 ( .A1(G234), .A2(n595), .ZN(n485) );
  XNOR2_X1 U582 ( .A(KEYINPUT20), .B(n485), .ZN(n488) );
  NAND2_X1 U583 ( .A1(n488), .A2(G217), .ZN(n486) );
  XOR2_X1 U584 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n490) );
  NAND2_X1 U585 ( .A1(n488), .A2(G221), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n490), .B(n489), .ZN(n633) );
  NAND2_X1 U587 ( .A1(G237), .A2(G234), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n491), .B(KEYINPUT14), .ZN(n631) );
  NOR2_X1 U589 ( .A1(G902), .A2(n714), .ZN(n493) );
  NOR2_X1 U590 ( .A1(G953), .A2(G952), .ZN(n492) );
  NOR2_X1 U591 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND2_X1 U592 ( .A1(G953), .A2(G900), .ZN(n495) );
  NAND2_X1 U593 ( .A1(n352), .A2(n495), .ZN(n531) );
  NOR2_X1 U594 ( .A1(n633), .A2(n531), .ZN(n496) );
  NAND2_X1 U595 ( .A1(n632), .A2(n496), .ZN(n535) );
  NOR2_X1 U596 ( .A1(n591), .A2(n535), .ZN(n497) );
  NAND2_X1 U597 ( .A1(n618), .A2(n497), .ZN(n498) );
  NAND2_X1 U598 ( .A1(G214), .A2(n525), .ZN(n647) );
  NAND2_X1 U599 ( .A1(n499), .A2(n647), .ZN(n550) );
  XOR2_X1 U600 ( .A(KEYINPUT110), .B(n550), .Z(n512) );
  XNOR2_X1 U601 ( .A(n500), .B(G107), .ZN(n515) );
  XNOR2_X1 U602 ( .A(n501), .B(n515), .ZN(n505) );
  NAND2_X1 U603 ( .A1(G227), .A2(n714), .ZN(n503) );
  XNOR2_X1 U604 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n508) );
  XNOR2_X2 U605 ( .A(n510), .B(n509), .ZN(n537) );
  XNOR2_X2 U606 ( .A(n537), .B(n511), .ZN(n635) );
  NAND2_X1 U607 ( .A1(n512), .A2(n635), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n514), .B(n513), .ZN(n528) );
  XOR2_X1 U609 ( .A(G122), .B(KEYINPUT16), .Z(n517) );
  NAND2_X1 U610 ( .A1(G224), .A2(n714), .ZN(n518) );
  XNOR2_X1 U611 ( .A(n519), .B(KEYINPUT17), .ZN(n521) );
  NAND2_X1 U612 ( .A1(G210), .A2(n525), .ZN(n527) );
  INV_X1 U613 ( .A(KEYINPUT95), .ZN(n526) );
  INV_X1 U614 ( .A(n558), .ZN(n551) );
  INV_X1 U615 ( .A(n647), .ZN(n529) );
  INV_X1 U616 ( .A(n537), .ZN(n530) );
  XNOR2_X1 U617 ( .A(n633), .B(KEYINPUT98), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n555), .A2(n539), .ZN(n625) );
  NOR2_X1 U619 ( .A1(n534), .A2(n625), .ZN(n630) );
  NOR2_X1 U620 ( .A1(n569), .A2(n535), .ZN(n536) );
  XNOR2_X1 U621 ( .A(n536), .B(KEYINPUT28), .ZN(n538) );
  NAND2_X1 U622 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U623 ( .A1(n349), .A2(n647), .ZN(n652) );
  INV_X1 U624 ( .A(n539), .ZN(n554) );
  OR2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n649) );
  NOR2_X1 U626 ( .A1(n652), .A2(n649), .ZN(n540) );
  NOR2_X1 U627 ( .A1(n544), .A2(n664), .ZN(n541) );
  XNOR2_X1 U628 ( .A(n541), .B(KEYINPUT42), .ZN(n722) );
  NAND2_X1 U629 ( .A1(n558), .A2(n647), .ZN(n543) );
  NOR2_X1 U630 ( .A1(n544), .A2(n565), .ZN(n619) );
  NAND2_X1 U631 ( .A1(KEYINPUT82), .A2(n651), .ZN(n545) );
  NAND2_X1 U632 ( .A1(n619), .A2(n545), .ZN(n546) );
  NAND2_X1 U633 ( .A1(n546), .A2(KEYINPUT47), .ZN(n549) );
  INV_X1 U634 ( .A(n619), .ZN(n614) );
  XOR2_X1 U635 ( .A(KEYINPUT83), .B(n651), .Z(n587) );
  NOR2_X1 U636 ( .A1(KEYINPUT47), .A2(n587), .ZN(n547) );
  AND2_X1 U637 ( .A1(n651), .A2(KEYINPUT47), .ZN(n548) );
  XNOR2_X1 U638 ( .A(KEYINPUT36), .B(n552), .ZN(n553) );
  INV_X1 U639 ( .A(n635), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n553), .A2(n570), .ZN(n629) );
  NAND2_X1 U641 ( .A1(n555), .A2(n554), .ZN(n578) );
  NOR2_X1 U642 ( .A1(n556), .A2(n578), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n346), .A2(n557), .ZN(n617) );
  XNOR2_X1 U644 ( .A(n617), .B(KEYINPUT84), .ZN(n559) );
  NAND2_X1 U645 ( .A1(n629), .A2(n559), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U647 ( .A1(n649), .A2(n564), .ZN(n568) );
  NAND2_X1 U648 ( .A1(G898), .A2(G953), .ZN(n566) );
  INV_X1 U649 ( .A(n569), .ZN(n640) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(KEYINPUT32), .Z(n572) );
  AND2_X1 U651 ( .A1(n570), .A2(n632), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n579), .A2(KEYINPUT44), .ZN(n573) );
  XNOR2_X1 U653 ( .A(n573), .B(KEYINPUT66), .ZN(n583) );
  XOR2_X1 U654 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n574) );
  XNOR2_X1 U655 ( .A(n576), .B(n575), .ZN(n663) );
  XNOR2_X1 U656 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n724), .A2(n579), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n724), .B(n580), .ZN(n581) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT31), .ZN(n624) );
  NAND2_X1 U660 ( .A1(n585), .A2(n356), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT100), .B(n586), .ZN(n607) );
  NAND2_X1 U662 ( .A1(n624), .A2(n607), .ZN(n589) );
  INV_X1 U663 ( .A(n587), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n632), .A2(n590), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n604) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT2), .ZN(n667) );
  NOR2_X2 U668 ( .A1(n667), .A2(n595), .ZN(n694) );
  NAND2_X1 U669 ( .A1(n694), .A2(G472), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT62), .B(KEYINPUT90), .Z(n596) );
  XNOR2_X1 U671 ( .A(n599), .B(n598), .ZN(n601) );
  NOR2_X1 U672 ( .A1(G952), .A2(n714), .ZN(n600) );
  XNOR2_X1 U673 ( .A(KEYINPUT92), .B(n600), .ZN(n693) );
  NAND2_X1 U674 ( .A1(n601), .A2(n698), .ZN(n603) );
  XOR2_X1 U675 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n602) );
  XNOR2_X1 U676 ( .A(n603), .B(n602), .ZN(G57) );
  XNOR2_X1 U677 ( .A(G101), .B(n604), .ZN(G3) );
  NOR2_X1 U678 ( .A1(n607), .A2(n622), .ZN(n605) );
  XOR2_X1 U679 ( .A(KEYINPUT114), .B(n605), .Z(n606) );
  XNOR2_X1 U680 ( .A(G104), .B(n606), .ZN(G6) );
  NOR2_X1 U681 ( .A1(n625), .A2(n607), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n609) );
  XNOR2_X1 U683 ( .A(G107), .B(KEYINPUT27), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n611), .B(n610), .ZN(G9) );
  XNOR2_X1 U686 ( .A(G110), .B(KEYINPUT116), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n613), .B(n612), .ZN(G12) );
  NOR2_X1 U688 ( .A1(n625), .A2(n614), .ZN(n616) );
  XNOR2_X1 U689 ( .A(G128), .B(KEYINPUT29), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(G30) );
  XNOR2_X1 U691 ( .A(G143), .B(n617), .ZN(G45) );
  XOR2_X1 U692 ( .A(G146), .B(KEYINPUT117), .Z(n621) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(G48) );
  NOR2_X1 U695 ( .A1(n622), .A2(n624), .ZN(n623) );
  XOR2_X1 U696 ( .A(G113), .B(n623), .Z(G15) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U698 ( .A(KEYINPUT118), .B(n626), .Z(n627) );
  XNOR2_X1 U699 ( .A(G116), .B(n627), .ZN(G18) );
  XOR2_X1 U700 ( .A(G125), .B(KEYINPUT37), .Z(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G27) );
  XOR2_X1 U702 ( .A(G134), .B(n630), .Z(G36) );
  NAND2_X1 U703 ( .A1(G952), .A2(n631), .ZN(n661) );
  XNOR2_X1 U704 ( .A(KEYINPUT121), .B(KEYINPUT52), .ZN(n659) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U706 ( .A(KEYINPUT49), .B(n634), .Z(n642) );
  NAND2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT119), .ZN(n638) );
  XNOR2_X1 U709 ( .A(KEYINPUT50), .B(n638), .ZN(n639) );
  NOR2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT51), .B(n645), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n664), .A2(n646), .ZN(n657) );
  NOR2_X1 U715 ( .A1(n349), .A2(n647), .ZN(n648) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT120), .ZN(n654) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n390), .A2(n655), .ZN(n656) );
  NOR2_X1 U721 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U722 ( .A(n659), .B(n658), .Z(n660) );
  NOR2_X1 U723 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U724 ( .A(n662), .B(KEYINPUT122), .ZN(n666) );
  NOR2_X1 U725 ( .A1(n664), .A2(n390), .ZN(n665) );
  NOR2_X1 U726 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U727 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U728 ( .A1(n669), .A2(G953), .ZN(n670) );
  XNOR2_X1 U729 ( .A(n670), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U730 ( .A(KEYINPUT56), .B(KEYINPUT86), .Z(n677) );
  NAND2_X1 U731 ( .A1(G210), .A2(n694), .ZN(n675) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT88), .ZN(n673) );
  XOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n672) );
  XNOR2_X1 U734 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n694), .A2(G469), .ZN(n681) );
  XOR2_X1 U736 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U737 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U738 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n693), .A2(n682), .ZN(G54) );
  NAND2_X1 U740 ( .A1(n694), .A2(G475), .ZN(n686) );
  XOR2_X1 U741 ( .A(KEYINPUT59), .B(KEYINPUT91), .Z(n683) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U743 ( .A1(n687), .A2(n698), .ZN(n689) );
  XOR2_X1 U744 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n688) );
  XNOR2_X1 U745 ( .A(n689), .B(n688), .ZN(G60) );
  NAND2_X1 U746 ( .A1(G478), .A2(n694), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(G63) );
  NAND2_X1 U749 ( .A1(G217), .A2(n694), .ZN(n697) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(n699) );
  INV_X1 U751 ( .A(G898), .ZN(n702) );
  NAND2_X1 U752 ( .A1(G953), .A2(G224), .ZN(n700) );
  XOR2_X1 U753 ( .A(KEYINPUT61), .B(n700), .Z(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n705) );
  NOR2_X1 U755 ( .A1(G953), .A2(n703), .ZN(n704) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U757 ( .A1(G898), .A2(n714), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U759 ( .A(n709), .B(n708), .Z(G69) );
  XNOR2_X1 U760 ( .A(n710), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U761 ( .A(n711), .B(n712), .ZN(n716) );
  XNOR2_X1 U762 ( .A(n716), .B(n713), .ZN(n715) );
  NAND2_X1 U763 ( .A1(n715), .A2(n714), .ZN(n720) );
  XNOR2_X1 U764 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n717), .A2(G900), .ZN(n718) );
  NAND2_X1 U766 ( .A1(G953), .A2(n718), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n720), .A2(n719), .ZN(G72) );
  XOR2_X1 U768 ( .A(G137), .B(KEYINPUT126), .Z(n721) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(G39) );
  XOR2_X1 U770 ( .A(G122), .B(KEYINPUT125), .Z(n723) );
  XNOR2_X1 U771 ( .A(n724), .B(n723), .ZN(G24) );
  XNOR2_X1 U772 ( .A(G140), .B(n725), .ZN(G42) );
  XNOR2_X1 U773 ( .A(n726), .B(G119), .ZN(G21) );
  XOR2_X1 U774 ( .A(G131), .B(n727), .Z(G33) );
endmodule

