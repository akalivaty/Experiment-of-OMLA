//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT69), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT70), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(new_n460), .B2(G125), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT71), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n468), .B(G2105), .C1(new_n472), .C2(new_n464), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n467), .B2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n460), .A2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n460), .A2(G124), .A3(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n484), .B1(KEYINPUT73), .B2(new_n488), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G102), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n470), .B2(new_n471), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n498), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n485), .B2(new_n486), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n492), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n508), .A2(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n509), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n520), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n514), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n514), .B1(new_n518), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n509), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n536), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n541), .A2(new_n514), .B1(new_n518), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n509), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT74), .Z(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  AND2_X1   g127(.A1(G53), .A2(G543), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n513), .A2(KEYINPUT75), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n510), .A2(new_n512), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(KEYINPUT9), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n515), .B2(new_n516), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n556), .A2(new_n557), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n513), .A2(G91), .A3(new_n517), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n559), .A2(new_n564), .A3(new_n566), .A4(new_n567), .ZN(G299));
  XNOR2_X1  g143(.A(new_n532), .B(KEYINPUT78), .ZN(G286));
  INV_X1    g144(.A(new_n518), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G87), .ZN(new_n571));
  INV_X1    g146(.A(new_n514), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n509), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n570), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n572), .A2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n514), .B1(new_n518), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT79), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n586), .A2(new_n509), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n513), .A2(G92), .A3(new_n517), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n591), .A2(new_n592), .B1(G54), .B2(new_n572), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n517), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n509), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(new_n597), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G321));
  XOR2_X1   g178(.A(G321), .B(KEYINPUT81), .Z(G284));
  NOR2_X1   g179(.A1(G299), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G286), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n609), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n476), .A2(G2104), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT83), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n476), .A2(G135), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n460), .A2(G2105), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n622), .B1(new_n623), .B2(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2096), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n620), .A2(new_n621), .A3(new_n629), .ZN(G156));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n636), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  OAI211_X1 g230(.A(new_n652), .B(new_n653), .C1(new_n651), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n648), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n628), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(G2100), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n664), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT20), .Z(new_n671));
  AOI211_X1 g246(.A(new_n669), .B(new_n671), .C1(new_n664), .C2(new_n668), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  INV_X1    g251(.A(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G32), .ZN(new_n681));
  NAND3_X1  g256(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT26), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n466), .A2(G105), .A3(G2104), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT95), .Z(new_n685));
  INV_X1    g260(.A(G129), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n624), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n683), .B(new_n687), .C1(G141), .C2(new_n476), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n681), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT27), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G5), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G171), .B2(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(G1961), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT96), .B1(new_n627), .B2(new_n680), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT31), .B(G11), .Z(new_n698));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n680), .B1(new_n699), .B2(G28), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT97), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n700), .A2(new_n701), .B1(new_n699), .B2(G28), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n680), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n692), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n692), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n691), .A2(new_n696), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(G164), .A2(new_n680), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G27), .B2(new_n680), .ZN(new_n714));
  INV_X1    g289(.A(G2078), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n692), .A2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n546), .B2(new_n692), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT89), .B(G1341), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n714), .A2(new_n715), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n712), .A2(new_n716), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT91), .B(KEYINPUT25), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G139), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n475), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n460), .A2(G127), .ZN(new_n730));
  NAND2_X1  g305(.A1(G115), .A2(G2104), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n466), .B2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G33), .B(new_n733), .S(G29), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n692), .A2(G4), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n602), .B2(new_n692), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1348), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n680), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n680), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n735), .B(new_n738), .C1(G2090), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G2090), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n737), .B2(G1348), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT24), .B(G34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(new_n680), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  INV_X1    g322(.A(G160), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n680), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n742), .A2(new_n744), .A3(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n734), .A2(G2072), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n680), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n476), .A2(G140), .ZN(new_n757));
  INV_X1    g332(.A(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n757), .B1(new_n758), .B2(new_n624), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n761), .A2(KEYINPUT90), .A3(G29), .ZN(new_n762));
  AOI21_X1  g337(.A(KEYINPUT90), .B1(new_n761), .B2(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2067), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n692), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G299), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n692), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n722), .A2(new_n752), .A3(new_n754), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G6), .B(G305), .S(G16), .Z(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G1981), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G1981), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n692), .A2(G23), .ZN(new_n777));
  INV_X1    g352(.A(G288), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n692), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT33), .B(G1976), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT88), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n692), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n692), .ZN(new_n784));
  INV_X1    g359(.A(G1971), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n775), .A2(new_n776), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n692), .A2(G24), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT86), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n791));
  NOR2_X1   g366(.A1(G290), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n692), .B1(G290), .B2(new_n791), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G1986), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n680), .A2(G25), .ZN(new_n798));
  NOR2_X1   g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT84), .Z(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G119), .ZN(new_n803));
  INV_X1    g378(.A(G131), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n803), .A2(new_n624), .B1(new_n475), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n798), .B1(new_n807), .B2(new_n680), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT85), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT35), .B(G1991), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n795), .A2(new_n796), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n797), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n788), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT36), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n788), .A2(new_n819), .A3(new_n815), .A4(new_n816), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n772), .B1(new_n818), .B2(new_n820), .ZN(G311));
  XNOR2_X1  g396(.A(G311), .B(KEYINPUT98), .ZN(G150));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n595), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n509), .B1(new_n825), .B2(KEYINPUT99), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(KEYINPUT99), .B2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n572), .A2(G55), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n570), .A2(G93), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n546), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n601), .A2(new_n609), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT100), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n830), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n733), .B(new_n761), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n502), .A2(new_n503), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n490), .B2(new_n491), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n688), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n843), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(new_n466), .B2(G118), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n624), .A2(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n476), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n617), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n807), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n847), .A2(new_n854), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n627), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT101), .B1(new_n847), .B2(new_n854), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n855), .B(new_n860), .C1(new_n862), .C2(new_n856), .ZN(new_n863));
  OAI221_X1 g438(.A(new_n842), .B1(new_n857), .B2(new_n860), .C1(new_n861), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g440(.A(G868), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n830), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G303), .B(G288), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G290), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G305), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n870), .A2(G305), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n870), .A2(G305), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n868), .A3(new_n871), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n874), .A2(KEYINPUT103), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT103), .B1(new_n874), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n876), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(KEYINPUT42), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n602), .A2(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n601), .A2(new_n768), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n601), .A2(KEYINPUT102), .A3(new_n768), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n884), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n890), .B2(KEYINPUT41), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n831), .B(new_n612), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n887), .A2(new_n888), .B1(new_n768), .B2(new_n601), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n892), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n882), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n867), .B1(new_n896), .B2(new_n866), .ZN(G295));
  OAI21_X1  g472(.A(new_n867), .B1(new_n896), .B2(new_n866), .ZN(G331));
  NAND2_X1  g473(.A1(G301), .A2(new_n532), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(G286), .B2(G301), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(new_n831), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n831), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n885), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n894), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n907), .C1(new_n877), .C2(new_n878), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n891), .A2(new_n903), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n894), .B1(new_n902), .B2(new_n901), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n879), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n908), .A2(new_n912), .A3(new_n913), .A4(new_n842), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n842), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n891), .B2(new_n903), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(new_n879), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n918), .B2(new_n879), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n913), .A4(new_n908), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n916), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT43), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n921), .A2(KEYINPUT43), .A3(new_n908), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(G397));
  INV_X1    g505(.A(new_n844), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n492), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G160), .A2(G40), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(KEYINPUT106), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n796), .A3(new_n870), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT126), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n688), .B(G1996), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n761), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n806), .B(new_n811), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n947), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n942), .A2(KEYINPUT46), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT46), .B1(new_n942), .B2(new_n955), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n941), .B1(new_n688), .B2(new_n950), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  NAND2_X1  g535(.A1(new_n807), .A2(new_n810), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n951), .A2(new_n961), .B1(G2067), .B2(new_n761), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n942), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n954), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n778), .A2(G1976), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n966), .B(new_n463), .C1(new_n467), .C2(new_n473), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n845), .A2(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n965), .A2(new_n969), .A3(G8), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n578), .A2(new_n579), .A3(new_n677), .A4(new_n580), .ZN(new_n972));
  INV_X1    g547(.A(G48), .ZN(new_n973));
  INV_X1    g548(.A(G86), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n973), .A2(new_n514), .B1(new_n518), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(G1981), .B1(new_n975), .B2(new_n577), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT49), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n972), .B(new_n976), .C1(new_n978), .C2(KEYINPUT49), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(G8), .A3(new_n981), .A4(new_n969), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n965), .A2(new_n969), .A3(G8), .A4(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n971), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G303), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(new_n967), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n506), .A2(new_n933), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n935), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n968), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n967), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2090), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n990), .B(G8), .C1(new_n995), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n969), .A2(G8), .ZN(new_n1002));
  INV_X1    g577(.A(new_n972), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G288), .A2(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n982), .B2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n987), .A2(new_n1001), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n986), .A2(new_n1001), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n992), .A2(new_n994), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n785), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n967), .C1(KEYINPUT50), .C2(new_n993), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n990), .B1(new_n1013), .B2(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1007), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n996), .A2(new_n750), .A3(new_n998), .A4(new_n967), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n845), .B2(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(G40), .A3(G160), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n935), .A2(G1384), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n506), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n506), .B2(new_n1021), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1016), .B1(new_n1024), .B2(G1966), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(G8), .A3(new_n606), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1026), .A2(KEYINPUT110), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1007), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n995), .B2(new_n1000), .ZN(new_n1033));
  INV_X1    g608(.A(new_n990), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1032), .B(new_n1035), .C1(new_n1028), .C2(new_n1027), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1006), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(KEYINPUT111), .A2(KEYINPUT57), .ZN(new_n1038));
  NAND2_X1  g613(.A1(KEYINPUT111), .A2(KEYINPUT57), .ZN(new_n1039));
  AND3_X1   g614(.A1(G299), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(G299), .B2(new_n1039), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1011), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n994), .A2(new_n967), .A3(new_n991), .A4(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1348), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n937), .A2(new_n934), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n999), .A2(new_n1052), .B1(new_n1053), .B2(new_n949), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n601), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1044), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1044), .A2(new_n1042), .A3(KEYINPUT112), .A4(new_n1046), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1051), .A2(new_n1056), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n999), .A2(new_n1052), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n949), .ZN(new_n1063));
  AND4_X1   g638(.A1(KEYINPUT60), .A2(new_n1062), .A3(new_n601), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n601), .B1(new_n1054), .B2(KEYINPUT60), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1064), .A2(new_n1065), .B1(KEYINPUT60), .B2(new_n1054), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1047), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(KEYINPUT61), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1057), .A2(KEYINPUT61), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1049), .A2(new_n1069), .A3(new_n1050), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1049), .A2(new_n1069), .A3(KEYINPUT118), .A4(new_n1050), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n955), .A2(new_n994), .A3(new_n967), .A4(new_n991), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  AND2_X1   g651(.A1(new_n969), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1075), .A2(new_n1077), .A3(KEYINPUT115), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n992), .A2(new_n955), .A3(new_n994), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n969), .A2(new_n1076), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n546), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT116), .B1(new_n1083), .B2(KEYINPUT59), .ZN(new_n1084));
  INV_X1    g659(.A(new_n546), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT115), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n546), .C1(new_n1078), .C2(new_n1082), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT117), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1084), .A2(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1061), .B1(new_n1074), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n999), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n506), .A2(new_n1021), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT109), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n506), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1100), .A2(new_n967), .A3(new_n1018), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n715), .A2(KEYINPUT53), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1098), .A2(G1961), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n994), .A2(new_n715), .A3(new_n991), .A4(new_n967), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1104), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n1112), .B2(G301), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1103), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1024), .A2(new_n1114), .B1(new_n999), .B2(new_n695), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1111), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(G171), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1098), .A2(G1961), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n465), .A2(new_n466), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n715), .A2(KEYINPUT123), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n715), .A2(KEYINPUT123), .ZN(new_n1123));
  OAI211_X1 g698(.A(KEYINPUT53), .B(G40), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1121), .A2(new_n463), .A3(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n936), .A2(new_n991), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1120), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(G301), .C1(new_n1109), .C2(new_n1116), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1113), .A2(new_n1119), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1025), .B2(new_n532), .ZN(new_n1133));
  OAI211_X1 g708(.A(G168), .B(new_n1016), .C1(new_n1024), .C2(G1966), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G8), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1132), .B1(new_n1134), .B2(G8), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT119), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1102), .A2(new_n710), .ZN(new_n1139));
  AOI21_X1  g714(.A(G168), .B1(new_n1139), .B2(new_n1016), .ZN(new_n1140));
  OAI211_X1 g715(.A(G8), .B(new_n1134), .C1(new_n1140), .C2(new_n1132), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(KEYINPUT51), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1112), .A2(G301), .ZN(new_n1146));
  AOI211_X1 g721(.A(new_n1126), .B(new_n1120), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1146), .B(KEYINPUT54), .C1(new_n1147), .C2(G301), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1131), .A2(new_n1145), .A3(new_n1015), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1037), .B1(new_n1097), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1119), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1118), .B1(new_n1117), .B2(G171), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1015), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1143), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1145), .B2(KEYINPUT62), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT124), .B(new_n1157), .C1(new_n1138), .C2(new_n1144), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT125), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1158), .B(new_n1164), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1150), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n942), .A2(G1986), .A3(G290), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n1167), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT107), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n953), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n964), .B1(new_n1166), .B2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g746(.A1(new_n661), .A2(G319), .A3(new_n646), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G229), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n923), .A2(new_n1174), .A3(new_n864), .ZN(G225));
  INV_X1    g749(.A(G225), .ZN(G308));
endmodule


