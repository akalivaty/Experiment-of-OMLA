//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT65), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G136), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OR2_X1    g056(.A1(G102), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G2105), .B1(KEYINPUT66), .B2(G114), .ZN(new_n483));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G114), .ZN(new_n484));
  OAI211_X1 g059(.A(G2104), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n486), .C2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT67), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n458), .C1(new_n486), .C2(new_n469), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n461), .A2(new_n494), .A3(G138), .A4(new_n458), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n490), .A2(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  AND2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(G50), .A3(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n498), .A2(new_n497), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n502), .A2(new_n510), .ZN(G166));
  NOR2_X1   g086(.A1(new_n497), .A2(new_n498), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT69), .B(G51), .Z(new_n515));
  AND2_X1   g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(new_n515), .B1(new_n503), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT7), .Z(new_n522));
  INV_X1    g097(.A(new_n509), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n522), .B1(G89), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n519), .A2(new_n520), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G168));
  NAND2_X1  g101(.A1(new_n514), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n509), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n505), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  OR3_X1    g107(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n529), .B2(new_n531), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n514), .A2(G43), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n509), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n505), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(G188));
  AOI22_X1  g121(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n505), .ZN(new_n548));
  OAI211_X1 g123(.A(G53), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n503), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n509), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n553), .A3(G91), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(G299));
  INV_X1    g130(.A(G171), .ZN(G301));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n525), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT73), .A4(new_n520), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  NAND3_X1  g137(.A1(new_n551), .A2(new_n553), .A3(G87), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n507), .A2(new_n508), .ZN(new_n564));
  INV_X1    g139(.A(G74), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G49), .A2(new_n514), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT74), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  AND3_X1   g145(.A1(KEYINPUT75), .A2(G73), .A3(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(G73), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n507), .B2(new_n508), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n505), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(KEYINPUT76), .B1(G48), .B2(new_n514), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n505), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n551), .A2(new_n553), .A3(G86), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n514), .A2(G47), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n509), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n505), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n564), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n514), .B2(G54), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n551), .A2(new_n553), .A3(G92), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  MUX2_X1   g175(.A(new_n600), .B(G301), .S(G868), .Z(G321));
  XNOR2_X1  g176(.A(G321), .B(KEYINPUT77), .ZN(G284));
  NOR2_X1   g177(.A1(G299), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n560), .B2(G868), .ZN(G297));
  AOI21_X1  g179(.A(new_n603), .B1(new_n560), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT78), .Z(G148));
  NAND2_X1  g183(.A1(new_n599), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g187(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n613));
  INV_X1    g188(.A(G111), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G2105), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n473), .A2(G135), .ZN(new_n616));
  AOI211_X1 g191(.A(new_n615), .B(new_n616), .C1(G123), .C2(new_n478), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT79), .B(G2096), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n461), .A2(new_n459), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2100), .Z(new_n623));
  NOR2_X1   g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(G156));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n629), .B(new_n635), .Z(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT17), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n642), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(new_n645), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g225(.A1(new_n644), .A2(new_n645), .B1(new_n650), .B2(KEYINPUT81), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(KEYINPUT81), .B2(new_n650), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT82), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n648), .A2(new_n646), .A3(new_n645), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  OR2_X1    g230(.A1(new_n647), .A2(new_n645), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n655), .C1(new_n644), .C2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2096), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n661), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n661), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT83), .B(KEYINPUT84), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G229));
  INV_X1    g256(.A(G29), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G26), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n473), .A2(G140), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT94), .ZN(new_n686));
  OR2_X1    g261(.A1(G104), .A2(G2105), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n687), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT95), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G128), .B2(new_n478), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n684), .B1(new_n692), .B2(new_n682), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT96), .B(G2067), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G16), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G5), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(G171), .B2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(G20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT23), .ZN(new_n702));
  INV_X1    g277(.A(G299), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n696), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1956), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n682), .A2(G35), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G162), .B2(new_n682), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT29), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n700), .B(new_n705), .C1(G2090), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G4), .A2(G16), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n599), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT91), .B(G1348), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n711), .B(new_n712), .Z(new_n713));
  NOR3_X1   g288(.A1(new_n695), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n696), .A2(G19), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n541), .B2(new_n696), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT92), .B(G1341), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n708), .A2(G2090), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G164), .A2(new_n682), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G27), .B2(new_n682), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n473), .A2(G141), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n459), .A2(G105), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT26), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n727), .B(new_n729), .C1(G129), .C2(new_n478), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G29), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n732), .B(KEYINPUT97), .C1(G29), .C2(G32), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(KEYINPUT97), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT27), .B(G1996), .Z(new_n735));
  OAI21_X1  g310(.A(new_n725), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n617), .A2(G29), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n682), .B1(new_n738), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n738), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G160), .B2(G29), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G2084), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n744), .A2(new_n682), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n737), .A2(new_n742), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n682), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n458), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n473), .B2(G139), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n682), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2072), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n721), .A2(new_n736), .A3(new_n748), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n696), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n696), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT98), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n759), .A2(G1966), .B1(new_n723), .B2(new_n724), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n734), .B2(new_n735), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n714), .A2(new_n757), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT99), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n696), .A2(G6), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n581), .B2(new_n696), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT32), .B(G1981), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT89), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n768), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n696), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n696), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1971), .ZN(new_n775));
  MUX2_X1   g350(.A(G23), .B(new_n568), .S(G16), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT33), .B(G1976), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n771), .A2(new_n772), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(KEYINPUT34), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G25), .A2(G29), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n473), .A2(G131), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n478), .A2(G119), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT86), .ZN(new_n786));
  INV_X1    g361(.A(G95), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n787), .A2(new_n458), .A3(KEYINPUT87), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT87), .B1(new_n787), .B2(new_n458), .ZN(new_n789));
  OAI221_X1 g364(.A(G2104), .B1(G107), .B2(new_n458), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n784), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n783), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT35), .B(G1991), .Z(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n696), .A2(G24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n588), .B2(new_n696), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1986), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n796), .B(new_n801), .C1(new_n780), .C2(KEYINPUT34), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n782), .A2(new_n802), .A3(KEYINPUT90), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT90), .B1(new_n782), .B2(new_n802), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n803), .A2(KEYINPUT36), .A3(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(KEYINPUT36), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n765), .A2(new_n805), .A3(new_n806), .ZN(G150));
  INV_X1    g382(.A(G150), .ZN(G311));
  NAND2_X1  g383(.A1(new_n599), .A2(G559), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT38), .Z(new_n810));
  AOI22_X1  g385(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(new_n505), .ZN(new_n812));
  AOI22_X1  g387(.A1(G93), .A2(new_n523), .B1(new_n514), .B2(G55), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n541), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n810), .B(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n814), .A2(new_n818), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n791), .B(new_n621), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n473), .A2(G142), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n458), .A2(G118), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT101), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n826), .B2(KEYINPUT101), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n827), .A2(new_n829), .B1(new_n478), .B2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n824), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n493), .A2(new_n495), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n485), .A2(new_n487), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n832), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n691), .B(new_n754), .ZN(new_n837));
  INV_X1    g412(.A(new_n731), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(G160), .B(KEYINPUT100), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n480), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(new_n617), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n840), .A2(new_n848), .A3(new_n841), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g426(.A(G166), .B(KEYINPUT103), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n581), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n588), .B(new_n568), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n581), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n854), .B1(new_n853), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT42), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n815), .B(new_n609), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n599), .B(new_n703), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(KEYINPUT41), .B2(new_n861), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n862), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n859), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(G868), .B2(new_n814), .ZN(G295));
  OAI21_X1  g445(.A(new_n869), .B1(G868), .B2(new_n814), .ZN(G331));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n558), .A2(new_n559), .B1(new_n533), .B2(new_n534), .ZN(new_n873));
  NOR2_X1   g448(.A1(G171), .A2(G168), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n815), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n560), .A2(G171), .ZN(new_n877));
  INV_X1    g452(.A(new_n815), .ZN(new_n878));
  NAND2_X1  g453(.A1(G301), .A2(new_n525), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  MUX2_X1   g457(.A(new_n863), .B(KEYINPUT41), .S(new_n861), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n861), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n875), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n858), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n876), .A2(new_n886), .A3(new_n881), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n880), .A2(new_n875), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n866), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n866), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n858), .B(new_n891), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n890), .A2(KEYINPUT106), .A3(new_n896), .A4(new_n847), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n847), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n858), .B1(new_n884), .B2(new_n887), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n872), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n889), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT43), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n872), .B1(new_n903), .B2(new_n905), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT43), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(G397));
  INV_X1    g487(.A(KEYINPUT127), .ZN(new_n913));
  AOI21_X1  g488(.A(G1384), .B1(new_n833), .B2(new_n834), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n914), .B2(KEYINPUT107), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G40), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n464), .A2(new_n467), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1996), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n921), .A2(new_n922), .A3(new_n731), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT109), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n691), .B(G2067), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n838), .A2(G1996), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G1986), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n588), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT108), .Z(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n931), .B2(new_n588), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n925), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n791), .B(new_n795), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n925), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n490), .A2(new_n491), .ZN(new_n939));
  AOI21_X1  g514(.A(G1384), .B1(new_n939), .B2(new_n833), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT50), .B(G1384), .C1(new_n833), .C2(new_n834), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n940), .A2(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G2084), .ZN(new_n945));
  OAI211_X1 g520(.A(KEYINPUT110), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n920), .A4(new_n946), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n459), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n465), .A2(new_n466), .ZN(new_n949));
  OAI211_X1 g524(.A(G40), .B(new_n948), .C1(new_n949), .C2(new_n458), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n835), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n952), .B2(new_n916), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n485), .A2(KEYINPUT67), .A3(new_n487), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT67), .B1(new_n485), .B2(new_n487), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n833), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1966), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n947), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G8), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n962), .A2(G286), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(G166), .B2(new_n965), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT55), .B(G8), .C1(new_n502), .C2(new_n510), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1971), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n835), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n920), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT45), .B1(new_n956), .B2(new_n951), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n956), .A2(new_n941), .A3(new_n951), .ZN(new_n974));
  INV_X1    g549(.A(G2090), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n488), .B1(new_n493), .B2(new_n495), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT50), .B1(new_n976), .B2(G1384), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(new_n920), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n968), .B1(new_n979), .B2(G8), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n963), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n941), .B1(new_n956), .B2(new_n951), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n943), .B1(new_n914), .B2(new_n941), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n946), .B(new_n920), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n985), .B2(G2090), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(G8), .A3(new_n968), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n986), .A2(KEYINPUT111), .A3(G8), .A4(new_n968), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n965), .B1(new_n920), .B2(new_n914), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n568), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT52), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n569), .B2(G1976), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  OAI211_X1 g574(.A(G48), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n1000));
  INV_X1    g575(.A(G86), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n509), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(G1981), .B1(new_n1002), .B2(new_n575), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT112), .B(G1981), .C1(new_n1002), .C2(new_n575), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1981), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n576), .A2(new_n579), .A3(new_n1008), .A4(new_n580), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT49), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n993), .B(new_n1010), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n581), .A2(new_n1008), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1014), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n1010), .A2(new_n993), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT113), .B1(new_n1014), .B2(KEYINPUT49), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n999), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n992), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g598(.A(G1976), .B(G288), .C1(new_n1016), .C2(new_n1021), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1009), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n993), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n963), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n968), .B1(new_n986), .B2(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT63), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1023), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n999), .B(new_n980), .C1(new_n1016), .C2(new_n1021), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n991), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1031), .B2(new_n991), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n971), .A2(new_n972), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n724), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1035), .A2(new_n1037), .B1(new_n985), .B2(new_n699), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT124), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n958), .B2(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n724), .A4(new_n957), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G171), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n533), .A2(KEYINPUT54), .A3(new_n534), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n918), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT125), .B(G2078), .Z(new_n1049));
  NOR3_X1   g624(.A1(new_n971), .A2(new_n1035), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1047), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1043), .A2(new_n1047), .B1(new_n1051), .B2(new_n1038), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(G8), .C1(new_n961), .C2(new_n525), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n525), .A2(G8), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT123), .B1(new_n961), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1058), .B(new_n1055), .C1(new_n947), .C2(new_n960), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1054), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1053), .B(new_n1056), .C1(new_n961), .C2(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1052), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1033), .A2(new_n1034), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n985), .A2(new_n712), .ZN(new_n1064));
  INV_X1    g639(.A(G2067), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n920), .A2(new_n1065), .A3(new_n914), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT118), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT60), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n599), .B2(KEYINPUT121), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n599), .A2(KEYINPUT121), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1064), .A2(new_n1067), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1064), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1070), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT60), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n550), .B2(KEYINPUT116), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(G299), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n972), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n950), .B1(KEYINPUT45), .B2(new_n914), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(G2072), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT115), .B(G1956), .Z(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n950), .B1(new_n952), .B2(KEYINPUT50), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n974), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1082), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n974), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n977), .A2(new_n920), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1081), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(new_n1098), .A3(KEYINPUT61), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(new_n1096), .A3(new_n1081), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1079), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1104), .B2(new_n1082), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT120), .A4(new_n1098), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n1071), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT58), .B(G1341), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n920), .B2(new_n914), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1036), .B2(new_n922), .ZN(new_n1113));
  INV_X1    g688(.A(new_n541), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1113), .A2(KEYINPUT59), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT59), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1078), .A2(new_n1108), .A3(new_n1109), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1092), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n600), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1100), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1030), .B1(new_n1063), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1031), .A2(new_n991), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT126), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1043), .A2(G171), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n962), .A2(KEYINPUT51), .A3(new_n1055), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1054), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1126), .B1(new_n1128), .B2(KEYINPUT62), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1060), .A2(KEYINPUT62), .A3(new_n1061), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1031), .A2(new_n1032), .A3(new_n991), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n938), .B1(new_n1123), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n925), .A2(new_n922), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT46), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n925), .B1(new_n926), .B2(new_n838), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT47), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n792), .A2(new_n794), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n929), .A2(new_n1139), .B1(G2067), .B2(new_n691), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n925), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n933), .A2(new_n921), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT48), .Z(new_n1143));
  NAND3_X1  g718(.A1(new_n930), .A2(new_n937), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n913), .B1(new_n1133), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1030), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1125), .A2(new_n1131), .A3(new_n1128), .A4(new_n1052), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(new_n1132), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n938), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1145), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT127), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1146), .A2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g730(.A(G319), .B1(new_n639), .B2(new_n640), .ZN(new_n1157));
  NOR2_X1   g731(.A1(G227), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n850), .A2(new_n680), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g733(.A1(new_n909), .A2(new_n910), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n1159), .A2(new_n1160), .ZN(G308));
  OR2_X1    g735(.A1(new_n1159), .A2(new_n1160), .ZN(G225));
endmodule


