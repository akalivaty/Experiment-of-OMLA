

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(G543), .B(KEYINPUT0), .Z(n520) );
  AND2_X1 U555 ( .A1(G1976), .A2(G288), .ZN(n521) );
  OR2_X1 U556 ( .A1(n723), .A2(n717), .ZN(n522) );
  NOR2_X1 U557 ( .A1(n723), .A2(n521), .ZN(n523) );
  AND2_X1 U558 ( .A1(n715), .A2(n523), .ZN(n524) );
  XOR2_X1 U559 ( .A(KEYINPUT31), .B(n693), .Z(n525) );
  AND2_X1 U560 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U561 ( .A(n713), .B(KEYINPUT100), .ZN(n721) );
  NAND2_X1 U562 ( .A1(n938), .A2(n522), .ZN(n718) );
  OR2_X1 U563 ( .A1(n719), .A2(n718), .ZN(n726) );
  XNOR2_X1 U564 ( .A(n530), .B(n529), .ZN(n882) );
  XNOR2_X1 U565 ( .A(KEYINPUT15), .B(n653), .ZN(n900) );
  NOR2_X1 U566 ( .A1(G651), .A2(n586), .ZN(n782) );
  NOR2_X1 U567 ( .A1(n544), .A2(n543), .ZN(G160) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U569 ( .A1(n885), .A2(G114), .ZN(n526) );
  XNOR2_X1 U570 ( .A(n526), .B(KEYINPUT88), .ZN(n528) );
  INV_X1 U571 ( .A(G2105), .ZN(n531) );
  AND2_X4 U572 ( .A1(n531), .A2(G2104), .ZN(n881) );
  NAND2_X1 U573 ( .A1(G102), .A2(n881), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n535) );
  XNOR2_X1 U575 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n530) );
  NOR2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G138), .A2(n882), .ZN(n533) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n531), .ZN(n886) );
  NAND2_X1 U579 ( .A1(G126), .A2(n886), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U581 ( .A1(n535), .A2(n534), .ZN(G164) );
  INV_X1 U582 ( .A(KEYINPUT23), .ZN(n537) );
  NAND2_X1 U583 ( .A1(G101), .A2(n881), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U585 ( .A(n538), .B(KEYINPUT64), .ZN(n540) );
  NAND2_X1 U586 ( .A1(G113), .A2(n885), .ZN(n539) );
  NAND2_X1 U587 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U588 ( .A1(G137), .A2(n882), .ZN(n542) );
  NAND2_X1 U589 ( .A1(G125), .A2(n886), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U591 ( .A(G651), .ZN(n549) );
  NOR2_X1 U592 ( .A1(G543), .A2(n549), .ZN(n546) );
  XNOR2_X1 U593 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n545) );
  XNOR2_X1 U594 ( .A(n546), .B(n545), .ZN(n778) );
  NAND2_X1 U595 ( .A1(G61), .A2(n778), .ZN(n548) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n779) );
  NAND2_X1 U597 ( .A1(G86), .A2(n779), .ZN(n547) );
  NAND2_X1 U598 ( .A1(n548), .A2(n547), .ZN(n552) );
  XNOR2_X1 U599 ( .A(KEYINPUT66), .B(n520), .ZN(n586) );
  NOR2_X1 U600 ( .A1(n549), .A2(n586), .ZN(n777) );
  NAND2_X1 U601 ( .A1(n777), .A2(G73), .ZN(n550) );
  XOR2_X1 U602 ( .A(KEYINPUT2), .B(n550), .Z(n551) );
  NOR2_X1 U603 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U604 ( .A1(n782), .A2(G48), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n554), .A2(n553), .ZN(G305) );
  NAND2_X1 U606 ( .A1(G64), .A2(n778), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G52), .A2(n782), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n561) );
  NAND2_X1 U609 ( .A1(G90), .A2(n779), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G77), .A2(n777), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n559), .Z(n560) );
  NOR2_X1 U613 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U614 ( .A1(n778), .A2(G63), .ZN(n562) );
  XNOR2_X1 U615 ( .A(n562), .B(KEYINPUT74), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G51), .A2(n782), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U618 ( .A(KEYINPUT6), .B(n565), .ZN(n572) );
  NAND2_X1 U619 ( .A1(n779), .A2(G89), .ZN(n566) );
  XNOR2_X1 U620 ( .A(n566), .B(KEYINPUT4), .ZN(n568) );
  NAND2_X1 U621 ( .A1(G76), .A2(n777), .ZN(n567) );
  NAND2_X1 U622 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U623 ( .A(KEYINPUT5), .B(n569), .ZN(n570) );
  XNOR2_X1 U624 ( .A(KEYINPUT73), .B(n570), .ZN(n571) );
  NOR2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(n573), .Z(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G75), .A2(n777), .ZN(n574) );
  XNOR2_X1 U629 ( .A(n574), .B(KEYINPUT84), .ZN(n577) );
  NAND2_X1 U630 ( .A1(G62), .A2(n778), .ZN(n575) );
  XOR2_X1 U631 ( .A(KEYINPUT83), .B(n575), .Z(n576) );
  NAND2_X1 U632 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U633 ( .A1(G88), .A2(n779), .ZN(n579) );
  NAND2_X1 U634 ( .A1(G50), .A2(n782), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U636 ( .A1(n581), .A2(n580), .ZN(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(G49), .A2(n782), .ZN(n583) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n582) );
  NAND2_X1 U640 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U641 ( .A1(n778), .A2(n584), .ZN(n585) );
  XNOR2_X1 U642 ( .A(n585), .B(KEYINPUT82), .ZN(n588) );
  NAND2_X1 U643 ( .A1(G87), .A2(n586), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n588), .A2(n587), .ZN(G288) );
  NAND2_X1 U645 ( .A1(G85), .A2(n779), .ZN(n590) );
  NAND2_X1 U646 ( .A1(G72), .A2(n777), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U648 ( .A1(G60), .A2(n778), .ZN(n592) );
  NAND2_X1 U649 ( .A1(G47), .A2(n782), .ZN(n591) );
  NAND2_X1 U650 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U651 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X1 U652 ( .A1(G164), .A2(G1384), .ZN(n626) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n624) );
  NOR2_X1 U654 ( .A1(n626), .A2(n624), .ZN(n744) );
  NAND2_X1 U655 ( .A1(G104), .A2(n881), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G140), .A2(n882), .ZN(n595) );
  NAND2_X1 U657 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U658 ( .A(KEYINPUT34), .B(n597), .Z(n604) );
  NAND2_X1 U659 ( .A1(n886), .A2(G128), .ZN(n598) );
  XOR2_X1 U660 ( .A(KEYINPUT89), .B(n598), .Z(n600) );
  NAND2_X1 U661 ( .A1(n885), .A2(G116), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U663 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n601) );
  XNOR2_X1 U664 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U665 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U666 ( .A(KEYINPUT36), .B(n605), .Z(n895) );
  XNOR2_X1 U667 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  OR2_X1 U668 ( .A1(n895), .A2(n742), .ZN(n606) );
  XNOR2_X1 U669 ( .A(n606), .B(KEYINPUT91), .ZN(n1013) );
  NAND2_X1 U670 ( .A1(n744), .A2(n1013), .ZN(n740) );
  XNOR2_X1 U671 ( .A(KEYINPUT92), .B(G1991), .ZN(n916) );
  NAND2_X1 U672 ( .A1(G107), .A2(n885), .ZN(n608) );
  NAND2_X1 U673 ( .A1(G95), .A2(n881), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U675 ( .A1(G131), .A2(n882), .ZN(n610) );
  NAND2_X1 U676 ( .A1(G119), .A2(n886), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n610), .A2(n609), .ZN(n611) );
  OR2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n892) );
  NAND2_X1 U679 ( .A1(n916), .A2(n892), .ZN(n621) );
  NAND2_X1 U680 ( .A1(G117), .A2(n885), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G129), .A2(n886), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n881), .A2(G105), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT38), .B(n615), .Z(n616) );
  NOR2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n882), .A2(G141), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n864) );
  NAND2_X1 U688 ( .A1(G1996), .A2(n864), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n995) );
  NAND2_X1 U690 ( .A1(n995), .A2(n744), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT93), .ZN(n736) );
  INV_X1 U692 ( .A(n736), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n740), .A2(n623), .ZN(n730) );
  INV_X1 U694 ( .A(n624), .ZN(n625) );
  NAND2_X2 U695 ( .A1(n626), .A2(n625), .ZN(n695) );
  NAND2_X1 U696 ( .A1(G8), .A2(n695), .ZN(n723) );
  NOR2_X1 U697 ( .A1(G1981), .A2(G305), .ZN(n627) );
  XOR2_X1 U698 ( .A(n627), .B(KEYINPUT24), .Z(n628) );
  NOR2_X1 U699 ( .A1(n723), .A2(n628), .ZN(n728) );
  INV_X1 U700 ( .A(n695), .ZN(n664) );
  NOR2_X1 U701 ( .A1(n664), .A2(G1961), .ZN(n632) );
  XOR2_X1 U702 ( .A(G2078), .B(KEYINPUT25), .Z(n922) );
  INV_X1 U703 ( .A(KEYINPUT94), .ZN(n629) );
  XNOR2_X2 U704 ( .A(n629), .B(n695), .ZN(n670) );
  INV_X1 U705 ( .A(n670), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n922), .A2(n630), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT95), .ZN(n686) );
  NAND2_X1 U709 ( .A1(n686), .A2(G171), .ZN(n685) );
  NAND2_X1 U710 ( .A1(G65), .A2(n778), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G53), .A2(n782), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G91), .A2(n779), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G78), .A2(n777), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n791) );
  NAND2_X1 U717 ( .A1(n670), .A2(G2072), .ZN(n641) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n641), .B(n640), .ZN(n643) );
  INV_X1 U720 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U721 ( .A1(n670), .A2(n969), .ZN(n642) );
  NOR2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n678) );
  OR2_X1 U723 ( .A1(n791), .A2(n678), .ZN(n644) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT28), .ZN(n682) );
  NAND2_X1 U725 ( .A1(G54), .A2(n782), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT72), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G66), .A2(n778), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G92), .A2(n779), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n777), .A2(G79), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT71), .ZN(n649) );
  NOR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U734 ( .A1(G56), .A2(n778), .ZN(n654) );
  XOR2_X1 U735 ( .A(KEYINPUT14), .B(n654), .Z(n661) );
  NAND2_X1 U736 ( .A1(G81), .A2(n779), .ZN(n655) );
  XOR2_X1 U737 ( .A(KEYINPUT12), .B(n655), .Z(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(KEYINPUT69), .ZN(n658) );
  NAND2_X1 U739 ( .A1(G68), .A2(n777), .ZN(n657) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U741 ( .A(KEYINPUT13), .B(n659), .Z(n660) );
  NOR2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n782), .A2(G43), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n954) );
  AND2_X1 U745 ( .A1(n664), .A2(G1996), .ZN(n666) );
  XNOR2_X1 U746 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n666), .B(n665), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n695), .A2(G1341), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U750 ( .A1(n954), .A2(n669), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n900), .A2(n675), .ZN(n674) );
  NAND2_X1 U752 ( .A1(G2067), .A2(n670), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G1348), .A2(n695), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n677) );
  OR2_X1 U756 ( .A1(n900), .A2(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n791), .A2(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U761 ( .A(KEYINPUT29), .B(n683), .Z(n684) );
  NAND2_X1 U762 ( .A1(n685), .A2(n684), .ZN(n694) );
  NOR2_X1 U763 ( .A1(G171), .A2(n686), .ZN(n687) );
  XNOR2_X1 U764 ( .A(n687), .B(KEYINPUT98), .ZN(n692) );
  NOR2_X1 U765 ( .A1(G1966), .A2(n723), .ZN(n708) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n695), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n708), .A2(n705), .ZN(n688) );
  NAND2_X1 U768 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U769 ( .A(KEYINPUT30), .B(n689), .ZN(n690) );
  NOR2_X1 U770 ( .A1(n690), .A2(G168), .ZN(n691) );
  NOR2_X1 U771 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U772 ( .A1(n694), .A2(n525), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n706), .A2(G286), .ZN(n702) );
  INV_X1 U774 ( .A(G8), .ZN(n700) );
  NOR2_X1 U775 ( .A1(G1971), .A2(n723), .ZN(n697) );
  NOR2_X1 U776 ( .A1(G2090), .A2(n695), .ZN(n696) );
  NOR2_X1 U777 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U778 ( .A1(n698), .A2(G303), .ZN(n699) );
  OR2_X1 U779 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U780 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n703) );
  XNOR2_X1 U781 ( .A(n704), .B(n703), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G8), .A2(n705), .ZN(n710) );
  INV_X1 U783 ( .A(n706), .ZN(n707) );
  NOR2_X1 U784 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U785 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U787 ( .A1(G1976), .A2(G288), .ZN(n716) );
  NOR2_X1 U788 ( .A1(G1971), .A2(G303), .ZN(n714) );
  NOR2_X1 U789 ( .A1(n716), .A2(n714), .ZN(n952) );
  NAND2_X1 U790 ( .A1(n721), .A2(n952), .ZN(n715) );
  NOR2_X1 U791 ( .A1(KEYINPUT33), .A2(n524), .ZN(n719) );
  XOR2_X1 U792 ( .A(G1981), .B(G305), .Z(n938) );
  NAND2_X1 U793 ( .A1(n716), .A2(KEYINPUT33), .ZN(n717) );
  NOR2_X1 U794 ( .A1(G2090), .A2(G303), .ZN(n720) );
  NAND2_X1 U795 ( .A1(G8), .A2(n720), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U798 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U801 ( .A(G1986), .B(G290), .ZN(n941) );
  NAND2_X1 U802 ( .A1(n941), .A2(n744), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n747) );
  NOR2_X1 U804 ( .A1(G1996), .A2(n864), .ZN(n992) );
  NOR2_X1 U805 ( .A1(n916), .A2(n892), .ZN(n998) );
  NOR2_X1 U806 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n998), .A2(n733), .ZN(n734) );
  XOR2_X1 U808 ( .A(KEYINPUT101), .B(n734), .Z(n735) );
  NOR2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U810 ( .A(n737), .B(KEYINPUT102), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n992), .A2(n738), .ZN(n739) );
  XNOR2_X1 U812 ( .A(KEYINPUT39), .B(n739), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n742), .A2(n895), .ZN(n1006) );
  NAND2_X1 U815 ( .A1(n743), .A2(n1006), .ZN(n745) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U818 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U819 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U820 ( .A1(G111), .A2(n885), .ZN(n750) );
  NAND2_X1 U821 ( .A1(G99), .A2(n881), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n756) );
  NAND2_X1 U823 ( .A1(n886), .A2(G123), .ZN(n751) );
  XNOR2_X1 U824 ( .A(n751), .B(KEYINPUT18), .ZN(n753) );
  NAND2_X1 U825 ( .A1(G135), .A2(n882), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U827 ( .A(KEYINPUT77), .B(n754), .Z(n755) );
  NOR2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U829 ( .A(KEYINPUT78), .B(n757), .Z(n1000) );
  XNOR2_X1 U830 ( .A(n1000), .B(G2096), .ZN(n758) );
  OR2_X1 U831 ( .A1(G2100), .A2(n758), .ZN(G156) );
  INV_X1 U832 ( .A(n791), .ZN(G299) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  INV_X1 U834 ( .A(G120), .ZN(G236) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n759) );
  XNOR2_X1 U838 ( .A(n759), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U839 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n761) );
  INV_X1 U840 ( .A(G223), .ZN(n814) );
  NAND2_X1 U841 ( .A1(G567), .A2(n814), .ZN(n760) );
  XNOR2_X1 U842 ( .A(n761), .B(n760), .ZN(G234) );
  INV_X1 U843 ( .A(n954), .ZN(n762) );
  NAND2_X1 U844 ( .A1(n762), .A2(G860), .ZN(G153) );
  INV_X1 U845 ( .A(G171), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G301), .A2(G868), .ZN(n763) );
  XNOR2_X1 U847 ( .A(n763), .B(KEYINPUT70), .ZN(n765) );
  INV_X1 U848 ( .A(G868), .ZN(n796) );
  INV_X1 U849 ( .A(n900), .ZN(n948) );
  NAND2_X1 U850 ( .A1(n796), .A2(n948), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(G284) );
  NOR2_X1 U852 ( .A1(G286), .A2(n796), .ZN(n767) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(G297) );
  INV_X1 U855 ( .A(G559), .ZN(n768) );
  NOR2_X1 U856 ( .A1(G860), .A2(n768), .ZN(n769) );
  XNOR2_X1 U857 ( .A(KEYINPUT75), .B(n769), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n770), .A2(n900), .ZN(n771) );
  XNOR2_X1 U859 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U860 ( .A1(G868), .A2(n954), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G868), .A2(n900), .ZN(n772) );
  NOR2_X1 U862 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U864 ( .A(KEYINPUT76), .B(n775), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G559), .A2(n900), .ZN(n776) );
  XOR2_X1 U866 ( .A(n954), .B(n776), .Z(n820) );
  NAND2_X1 U867 ( .A1(G80), .A2(n777), .ZN(n787) );
  NAND2_X1 U868 ( .A1(G67), .A2(n778), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G93), .A2(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n782), .A2(G55), .ZN(n783) );
  XOR2_X1 U872 ( .A(KEYINPUT80), .B(n783), .Z(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U875 ( .A(n788), .B(KEYINPUT81), .Z(n823) );
  XOR2_X1 U876 ( .A(n823), .B(G290), .Z(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(G305), .ZN(n790) );
  XOR2_X1 U878 ( .A(n790), .B(KEYINPUT19), .Z(n793) );
  XNOR2_X1 U879 ( .A(G166), .B(n791), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n794), .B(G288), .ZN(n899) );
  XNOR2_X1 U882 ( .A(n820), .B(n899), .ZN(n795) );
  NAND2_X1 U883 ( .A1(n795), .A2(G868), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n796), .A2(n823), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(G295) );
  NAND2_X1 U886 ( .A1(G2078), .A2(G2084), .ZN(n799) );
  XOR2_X1 U887 ( .A(KEYINPUT20), .B(n799), .Z(n800) );
  NAND2_X1 U888 ( .A1(G2090), .A2(n800), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT21), .B(n801), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n802), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U891 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U892 ( .A1(G220), .A2(G219), .ZN(n803) );
  XOR2_X1 U893 ( .A(KEYINPUT22), .B(n803), .Z(n804) );
  NOR2_X1 U894 ( .A1(G218), .A2(n804), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G96), .A2(n805), .ZN(n818) );
  NAND2_X1 U896 ( .A1(n818), .A2(G2106), .ZN(n811) );
  NOR2_X1 U897 ( .A1(G236), .A2(G237), .ZN(n806) );
  NAND2_X1 U898 ( .A1(G69), .A2(n806), .ZN(n807) );
  XNOR2_X1 U899 ( .A(KEYINPUT85), .B(n807), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n808), .A2(G108), .ZN(n809) );
  XNOR2_X1 U901 ( .A(KEYINPUT86), .B(n809), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n819), .A2(G567), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n911) );
  NAND2_X1 U904 ( .A1(G661), .A2(G483), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n911), .A2(n812), .ZN(n813) );
  XOR2_X1 U906 ( .A(KEYINPUT87), .B(n813), .Z(n817) );
  NAND2_X1 U907 ( .A1(n817), .A2(G36), .ZN(G176) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n814), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n815) );
  NAND2_X1 U910 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(G188) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(G325) );
  XNOR2_X1 U914 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U916 ( .A(G108), .ZN(G238) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U918 ( .A(KEYINPUT79), .B(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(G860), .A2(n821), .ZN(n822) );
  XOR2_X1 U920 ( .A(n823), .B(n822), .Z(G145) );
  XOR2_X1 U921 ( .A(G2454), .B(G2435), .Z(n825) );
  XNOR2_X1 U922 ( .A(G2438), .B(G2427), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n832) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(G2446), .Z(n827) );
  XNOR2_X1 U925 ( .A(G2443), .B(G2430), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U927 ( .A(n828), .B(G2451), .Z(n830) );
  XNOR2_X1 U928 ( .A(G1341), .B(G1348), .ZN(n829) );
  XNOR2_X1 U929 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n833), .A2(G14), .ZN(n834) );
  XOR2_X1 U932 ( .A(KEYINPUT104), .B(n834), .Z(G401) );
  XOR2_X1 U933 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U934 ( .A(G1996), .B(G1991), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n846) );
  XOR2_X1 U936 ( .A(KEYINPUT109), .B(G2474), .Z(n838) );
  XNOR2_X1 U937 ( .A(G1981), .B(KEYINPUT107), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(G1956), .B(G1961), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1966), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U943 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n846), .B(n845), .Z(G229) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2090), .B(KEYINPUT106), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n849), .B(G2678), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(G227) );
  NAND2_X1 U956 ( .A1(G124), .A2(n886), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n856), .B(KEYINPUT110), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G112), .A2(n885), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G100), .A2(n881), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G136), .A2(n882), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U964 ( .A1(n863), .A2(n862), .ZN(G162) );
  XNOR2_X1 U965 ( .A(n864), .B(G162), .ZN(n866) );
  XNOR2_X1 U966 ( .A(G164), .B(G160), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n880) );
  XOR2_X1 U968 ( .A(KEYINPUT113), .B(KEYINPUT112), .Z(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G118), .A2(n885), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G130), .A2(n886), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n881), .A2(G106), .ZN(n871) );
  XOR2_X1 U975 ( .A(KEYINPUT111), .B(n871), .Z(n873) );
  NAND2_X1 U976 ( .A1(n882), .A2(G142), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(n878), .B(n877), .Z(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n1002) );
  XNOR2_X1 U990 ( .A(n892), .B(n1002), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n1000), .B(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U994 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n954), .B(n899), .ZN(n902) );
  XNOR2_X1 U996 ( .A(G171), .B(n900), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n903), .B(G286), .ZN(n904) );
  NOR2_X1 U999 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(KEYINPUT114), .B(n905), .ZN(G397) );
  OR2_X1 U1001 ( .A1(n911), .A2(G401), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(n911), .ZN(G319) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1010 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n1016) );
  XOR2_X1 U1011 ( .A(G2090), .B(G35), .Z(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT119), .B(n912), .ZN(n928) );
  XNOR2_X1 U1013 ( .A(G2067), .B(G26), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G32), .B(G1996), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n921) );
  XOR2_X1 U1016 ( .A(G2072), .B(G33), .Z(n915) );
  NAND2_X1 U1017 ( .A1(n915), .A2(G28), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(KEYINPUT120), .B(n916), .ZN(n917) );
  XNOR2_X1 U1019 ( .A(G25), .B(n917), .ZN(n918) );
  NOR2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G27), .B(n922), .Z(n923) );
  XNOR2_X1 U1023 ( .A(KEYINPUT121), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT53), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT122), .ZN(n932) );
  XOR2_X1 U1028 ( .A(G2084), .B(G34), .Z(n930) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(n930), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n1016), .B(n933), .ZN(n935) );
  INV_X1 U1032 ( .A(G29), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(G11), .A2(n936), .ZN(n990) );
  INV_X1 U1035 ( .A(G16), .ZN(n986) );
  XNOR2_X1 U1036 ( .A(KEYINPUT56), .B(KEYINPUT123), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n986), .B(n937), .ZN(n960) );
  XNOR2_X1 U1038 ( .A(G1966), .B(G168), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n940), .B(KEYINPUT57), .ZN(n958) );
  NOR2_X1 U1041 ( .A1(n521), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(G1961), .B(G171), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(G1971), .A2(G303), .ZN(n942) );
  NAND2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(G1956), .B(G299), .ZN(n944) );
  NOR2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G1348), .B(n948), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n953), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1341), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n988) );
  XOR2_X1 U1056 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1060 ( .A(G1976), .B(KEYINPUT126), .Z(n963) );
  XNOR2_X1 U1061 ( .A(G23), .B(n963), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n967), .B(n966), .ZN(n983) );
  XNOR2_X1 U1064 ( .A(KEYINPUT125), .B(G1966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(n968), .B(G21), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G20), .B(n969), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1071 ( .A(KEYINPUT59), .B(G1348), .Z(n974) );
  XNOR2_X1 U1072 ( .A(G4), .B(n974), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(n977), .Z(n979) );
  XNOR2_X1 U1075 ( .A(G1961), .B(G5), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n984), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n1020) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT51), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1011) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT115), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT116), .B(n1001), .ZN(n1009) );
  XOR2_X1 U1092 ( .A(G2072), .B(n1002), .Z(n1004) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT50), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT117), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(G29), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

